��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� �����ޜ<(��l���R�l�iD�}�ŭ�L����6���8ﰘ~�Y�xI�h
�]�깵.�0i[�!:�N��~#<��3���~T���Ođ[/���e�fҾ����_6���*��"�������,TD�N�O'N��q��)����Q,�剺h�L�7R�*g�t�;�nG8T�����±m��d���}��٭;Z�����2���_���w��q��2�=��|׊U%|ggT��+� (`@ZĹ�KؚU�-)��w�)��,�g�A?�1�}��
̠��d�9���`ힸn%��Qq�a|S$���Z���	T�+���v?u&Q��xO3NXz�i�A��3A5o��k[U��jڊH w\�'�3�e�!�����(y�<�p�3N�.���ɴ����2_�c�H���[��#&n�D^�����E���&�$���5�7J��,��W�yk��p�}�/�9��z��l��}���S�����Gqz��ֺ� �쯺���h��^��SIm~ �����!V8=8�&1.�hn���Γ�-YК:�i�2�p	 �&7�ONz�M�?�ѕcДe��A���4�"�f�o�kG�~z��B���t�mU�.�u��j�wy�ѐ��eЧ�%\�Sg}��|��ѕ;)T`�������-��$��b����w�M����]��M�"��Ɣ�B!kuy��*T�Y*]�h������|�W-b}�kH��tw��y#�N��{A	�w	F���/���P��O���g��NE�r�e���_�n�'a��Id;�l���3��OUy��~���(�fct:E�\��ݭ[`ܶ��p޷�'G�Pq;�\�"������N)	"��KA~R�O���r�$�Ω=���r�gֱ��I���h� Pt}2��3WG��qT����ݡ�� �Iu2����nߖSFS����ᴬ�c�@Ϸ�Z	zY+�������w����W�q�9�u_U����4��T�æ�n�滠}�/��Jtž2ǎ㨔�2�^�qŀ�; �iq�w��M1h*��&��.��8x@�HUR��(��Ƚ�܍�=|=�Z�y�ɚVV��I��V/�����%�bb���{�J;��[hwWlX@�-S��XF@�l���������᎔�.e?�.Gi�u.�n[у�K�r27�A�nGL~�:%mp��%��O�������6��$۱O?d����LV���:\n*)���Y�=�|��ڗ��*O}�w9Gof�j���ox��tk��9�D�0�@8�~�&�<�TVpm*��e<]�Oem!żݺ�G���{+���_�;�,�[k&��h�#�S�:B��ߟ���}=��y�|9UV�;J�1v��?�\rQ��E<�ϙ�4!B�	0��Fg�f`��v�(N!�5�Z�zl�QUt�8[��~8�F�h��%����U �ڷ�R��������6Ǟ\�:�z������B�/IR,�T����o �e&�'������{��׽�!��q�%�L��J���*6ղ�BW�g�[�=�޷Baa��G�r�?[L(͛�ހ��"%m�b.�����k��!�t�>�7C�ص�ժ;�9��$����	�9\H4���0���b۫>ʠ_sMW���ٳ�(�U�`�b  7kej(��]�#�c�f����P�iA�,2�J{?���۔�jt\D#�o���C
rf�q!R�cc�3A��� y���-��O̊Yaג�T?#����}�*}�,�̙L0c�G��������v��Y�����"��zH�sb�tw�����%����W��bV�?x�b�,�g�M�/�?,v�6���U��&�����"�)̯�Ѓ�e�0
]ɻ^)WZ����jwV�(���E��ܺ	C�y�f��>���W��*� �����廬㣧��#
���VGz�JI�s?**��^�EǮ�p��N�vA~ ^��s3*��'��H��cmϭ@��H�+�JTo΁0�1���Y�	�Y��~�ב��i�6bybC�6��G��&3^�	C#q!�TTx����ӡ@������D�d@�]����`�3H����E�~9zl�"��3�a̭�^�𚧳�.*�^/�A<n� �V��L�IQ���=����^N8H�K�#$��)��l�S�^q/��W�.4%����`*9ܐ�UB����v��2]8��}d$[��g�ML�6�%���s�%�D�foCu[�.�����<ɗ/&�z�Z�o-/L���g����j
�3ц?���$R���6��K�~�=E~t<�	%�Ϳ���)��Z��}�QͰ���ޥ�ygWV�!�w���Xٷ��6'��%z/�7��Gy��w�X�n��Q�Ŏ��T�w�H1.0�� �=��7��2sGa3 )޳i�6�4�3�� �a�Q<7�����}0��̤]�k8TjR������ƶ��x���a�XŞ]!J��?���{xð�|�~ƶ��4���=�����d,�w]m�H&�-�>v��L�LK�L6�Lp=$�lB�jP<t<{��������E�Q�@���G�#��%�����Y���+63
P=�#�������Zj[b9ܒɶ�/�.��Җ;f�u:�zi�a����Ƨ?�j��i�2�ɓӗ����Ѡ����j��v?�t���t*a766��*N���}�KN+�S�@gO7Ks�4�\�㌝ѝܢ1�@sLj��jl�ɋjK���]A�3fi�]dou_l��nB��B�er�5�qf�����ɋ�
��@�CI���H�L�����\Hi:�o�����=�P�0��6)z��3�l�	�!���};���\�>��/��&b�T-*�~�����S������=�Q��|�-���u�� ���S6���L�N��KMܖ���7?�v
�_b&="�Μ����	82��U2?0��_���l�2��"��/ÜЦ0f��?d��:��}{�$��}io%�O=���F���0��L��D:�X�
�!}k2���n�$��ܭ��ٱPH�e���V���Mm�v=A�@��'��bKL�`F���P�ܗ|�	��i�@拗䎙ƙi4��)SVcVi�;���.�e ��궯��$��[�	9����O�]��S+-�6E4�Q�T��y��$<���`��7��o�2=Vm���qb���LD��'�	��q��D	�f�5�]cl{SC��Qf�-:��y�V�;��1���]�di�]^`#Lw�3�)��Ń�Na☟ Zo������!��MT�������'7(/^�Fp�X�X1�BW�7�E�h{�I�y�$�r�זa-ݺͷ}xlnțo%�.	�҉��iJ����u�6,̩h�Bz�_�M��1r	����z9�*�~�}�D%:�rF��ݘ�������L9��s�j�ۘ���v"��Ra#�Prj�$�$CUƤ����'|X�<�@��7m.�f�V5E��+�,����2�m�V�O�@����$�����ĝ�I+���f���t��H�l�Բ&�p�/���3Hw, j�u��;"l+�"�����X�s��`B��^�C)�������ƿ�����s���_}Lm-�\b��,E�+���IY��g�A���vCL���;�_��nK�0���$�i�[�X(�	����y!��y� ʸ���|=Fҡ�m�h*�����u��(���P]%*&e��sCwv���Ι�Fo�L�W���˕�o��$:��蛵y?Ԋ|�xF��r�M��Ft�
X.j�k��7#u�͍U�4ǎ�dM�\�#S�z����QA	���y�.��)���<E�u��:y���b�������T�M�R��d��A���:\�۩����pa��4������/qpU4	�7g#��Um��G��wV�Sjr5��:�J�Q��/i����n��TqYg���@��R�2Н��O�Rb�7�d�3wX��@Ol����u�dAl6�.S�
�]IN�`��s��e+jrr����{b�V별�d%���"���P{<�n������T,ǳx*�oX��f�r���8�\Ymc�T!;5����P����`�mB��FJ~_3$���9�RO��<�d;S���%��s�1�ܖ���c�%K��ݙ��x�N��1����q�Om��S��">CK�`�y�ȋ����A�����U@e����ş!^W��eZu�m� #y���,��f#U2O+Z �m�\fK�I���#Mk��0���Z+NDE,�.3���a�w�P���DLK4؁�7�ޓ�f(>��~�t��1��K�.���7���M:����b��a�{@q��N��
�ӕ�4�����G�����}��l`ӄ��W�&�F�򯕙�D��aw��o���N��]L�!McD�y�&:�V\$0�'��)S)�d[r�'5�����o4�hr�V��-��guT>��6!�-���j-�O�aw�6�Ȏ���Q������l�c��}�L}B�/�X�A�1Y_F�2��3���A��6U����^	��#��Q�1d;�����RNn$��YdUZ�K(���EnR��pV�)-��x^�~f:�'ym�;^�M�5��l�j�I3�8��އ-�6�eR�d M��L�P�E{P���Meδq��U�7G3 5���/���~�P{�vъS�,�_��7���t>�i�ۧ�D�L;�g����Z�Bn�%μ-v 6s�����ͅ2�8"�s�o�}�rY�I9n�� 	���W�.83/J2�,�M�T�{�?�Z@o��ڿ)���`����zQi|�w"��¿�f�}�w��#�൚ǽ)a���jl�zH��!��o�!���x<NJz�yR�?uR�6��fL�Dx�ߨS%�A�h//$��M�#�I�)���.���>L�#��a���R�%�v˭,W�ي����(���1���d�q�[��r������M0���a����Ƚ�g��!��N�O���w
W�)��9�"N� ���*���RM�"�բq��3z�d��s�l+n��TJ ��L3��k����_��*�xzaն��`�qJ��8p��䮚����{�#�/�2�0=8U�FD�<7��3�̖8���ҽ�H�b{��*�Ҷ�k�ٺ�0�i��;%0�z��7aA�%gĽCT&��F@�"6�_~N��$7�U5�bCxR��_f;���1g)%��+y��Lܛ��!��n�n �	�ц ��R�e ����Ho f-��)�?<7���LNP#X�-�=#ɹL���Ӏ)'ݳ�vd̋��"Xa��l��DN6|���e/���*�-�n�r6ϓe��Зg-�vPE�Д��)RSpR-Hd�2�w�џ�0EGs&jVX^�6�.�?�7�I�&���ߑd��v�%�]�s�X�_T���+Ly�e�>�_i�$9q����v�`�pS<v92�b���F��2�a.�����ɤ�R�/�� ��E�\ѷ�s*����DWPpe#�����	L��2��h%�I�V�w}�i�؋�#�!t�!_����^���5���D��L���m%��^����J����)���+C�J^�QPS�<-�S�	��N���O����́ӄ��7u�����.�ugP4	�5��y(�A���ZK��B�$ISd�-�NWJ�P&�.��>����nc�����B ���7���7;�-�����,����K��}u�0|���Mu��:!G�.��{u�5�]�6$zԃ}@��WB%�{9)�x
�4�l\��m�+�j9@sBCHӭ,�J�����_ CQO�_��&K�u�e���Q�E�H�Ըby������ 'U��{U�����E1'��CIhp��zʅ~4'.%�P�M��0��Q!|��\
n��^��o�s	�e�o(脴��p�xAӳ6 P�gAV���6��� wK��#v�>�:%���NR�l�-
9n9-��0��O�5~�)険��)�Kcs��/4��Ȥ�B5J�*����%�Am����J�fO�#�lG�Zs:��a<�vS��wP���LyIL|��Jx���ΎjTvJO�=��3��>�V!I�#qXn8}/8<����b9���2O�*zǭb��	�V�p��ૼfNK��ۨQl�K��lZtG�|9��:j˳v��%�r`����xT؁L��칈1`�^m�p�3�X	�FF>��n�L�/	[��7�.�ħ�=|�- t��ֵ�R�n�Y)��A�����Q�~�
��t9�K�ĩ����.y�m����M���]5����N�q:�r2xwsG3�ĝ!꒳E�	2 Z!�b�]*Y'�<R�Y�3��خ+�{�Z��:�)	{1�Wtj���Xnz�;��d��;Ē�;�S^�F`8@�Kh ��K�Q8����$��Y�Q�1)z�Ir�1{�U(g�WJ�;Q�m<����F���ۼ�$�U|�I�9���v�B�[k�QG���NO����2�ଢbX�j�A:hS�F�Kw�mo����4!� ���U���k8�z�y�7���=�K�[��-[M��Z��鹀F@�S�U���S��3U�߼���f����6�:|4�u�әG�����j�\�NA�Q��,���Lѯr�R�+t]ٰO�~k�����KU��E��z�K���`_ �܏���Hm�9����K¿�����c����Vr��٧���Nk:��F$�3�W�	%���U?g���؃19�4�Xphml���C��� #/:l�dW5S��O��9�%�;����V�0]�"`&}D	~D�"\���aIg�+ö�<�ۈ�pO�
<A1s)ŕo�F+���HUE�Z(0,4�ƿ��S K������M\ȕM�Ɍ���w˩�3�]&�$X��Y�͌f���,#����ڰ7C�u1h��E���iph�iL�YZ���F&&)'-	�}�#�����Pb������8[�΅��� �{�7ŠcP�p���o�mZ�M�7̮����M���_+x|��Q�/�j���n��#Å=�No�˭6o970�����!2�ƵB��|9A�Dט����5����0���RW��ljūQG:h@.�덒��ML>y�G��x'T8�l�ur�]�T�L? �!�@H�>S�8�,�E���{AmH_��o
K�:4�^���Tp�G�9"�{�T�y�tXb69 d��+i��	8��u6R�ZE/P�h���ILR�6��vg�����	�B�6��7��QX�܊)��2��I�KZ���ݗl�I�h_Bܔ���[.��ѿ�B%�:�Hh��4��Gp�/B*dÄ����]D��5����^�Teᘵ�?��Rؽ'nOO�F~O�M�rp2�J��Y'�Q&�oq���J���A~76ݓ���o�z��b�jPg�}��Q�_�Q*��<#�ڱ�b�H��Ӹ?�D;�Tg9���C/X�v�)4���!c�J
�M�vpF��E��`ㄍX;B�f�
]E��( ���:ӏ��.y��d�p�le�)��y��;�XN!�U4��%j�/<�����9�R�rd!n+F�<@u?�fu8�j��&�[r���L� �)�c$DV��6z�1��P��$Kt\j�Ja�;j]��G�ꎔ���܁��Hr
��|�����2�>b��1U�f̠4����#��]���4$���[�4���lj�@�JNJ��!{����m+C;��>�M�o.5`�b*As��y� ?����\�b�3f�E���Aӿ;�('1��h�S�ٺ�U�r���9�	}Pq�Lڛ?o��2U��Q<9Vb ���|D���
�j˿Ao���B����H3&���jD�7��/2;2�B�u�0��#���wނ�ބcb��F�eGA)�Ǩ���U.�֝>�
Hĵ���L�(~��3v&�P\�=j�<���,i�"_�6oJEf�"X�:��7*��K�f_rs��r�.?��I	^������.o��e�y��(k^'�B:Q����ڌ���f9�P�G��Hv�2��	:�L����8yQ���=@jw|�T=��a�O�PەBܴ��(�p\�!S���S�ےz~�ƽ5I���U��d�SE�n��i��\aά���Dx>w��y�l10�)�IÂ,	��Ų8T���'�]AJ�v�hYک���_!#u�u�p�M�#+"�*b{4��}��^�'
sL����ad�%��S���R@��!(���3O�����dI�[P�����@���K%����?�FBd:Z��j�B���q��m�na�6�L,���YO���a�-K���܋��3D5�Py@���^M�����rʓ<K���mC���׈&�u[��1L�ߢ���kW��:+�1��6p�5���M�H������g�u��R!��I=��u��m.�
�|��k7�)��fGt�J�������+�椟Xl�ųt��q%�(�Ng�(n#�B�g�M2��+��@H�2<{����6�[��G�j�v��3&)h���������O�Ϝ�܀��}`�2:���>s�S_[ù��+M��k�쁇���'��d�L���k����-F��Lp�t���|6�92L���:���'ȶ�97f�x�DQhT�D�ꉠ'.Rӫ��9Q�,|cp���L+��(td�:Q7&��Km,�}��&��(/�_D��
[��,�w� 
G.��7����ïv&n�J5�<�H"��s�(�&vJ�Iͬ�"д��s,������)T�h��?<HzC���\�����p��:���r��)OJoŶ�6��`�oXg����"��S=V�U.��q����ܷ<�B���p2+�|�g����5��/<�9+���#�oi���LC� (hh����葏�5hz�1�`���W#_{�\�B�)]�ic]��Ekb�ܽe�5o�l�&	��#�Br{\��4GF]�� u�  �94�6Aj��#�;f�e�/�L��*�w]��M\7`5�e��%'5h�`6`���N�=s�8(4�W�&5�k�#e$tᴦ���o�үM���N�H�G��Wn�H!e��ܱ��I��$�5/�x�L�ϴR�h��]D/�;�eX�'%G��8�n" `�ٔ+�"�=�JF����+:��|�|���uS��_e�C�C� �y��;�}�  d(=��I�)f<G�6k�<MB���XR�XW�m��1�g^ߝ����z�	/�a�!���z\bj�{"L:���Gl�����3�0���c1�g} V�wǘ��l7>��Q �V��t��n��Gk�U{#��!�j��/��[��k�W�*_�߶(��j��%	�0����
�v���_�3��Q1��-���Z�V�k�����Z�g�|W� �`8��Sqa9k�� �=D����6;/"��*����kVC۝�'U�QÅ���+����	�BO�����dd��W�v�=��y5�e*	)��tWE�:���1����?�gW+�`��8�-�u�n_Yh�L�9�9��������w� I���d��W�n�2�d&�
�RpRC�MPӞ�
wh�Yg,�`��$�vٱ��K���BY�����O�uc�}�L��g����c��"�l}f���G�Xe�-��{�5�My�Nr�F�e�}G��.+�м������n^M�%nٍ`�1أ�Q����9w�U�5��a��gs�fhǉ����re�r��z�k#dEG׌;=��������7�����T��{��&N��e��cGVL���\�:�aa:��F��?���Zzb&Zj*šW�����Һ�H��v��X��X`TV?KrL���}��cc�~��=�V�-D��B"�-�gFE�jF
AmUr�Y �~�
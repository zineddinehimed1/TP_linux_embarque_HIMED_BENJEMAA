��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"���99���{`���t���0�^���P���D�21�I�����Il:R4)dOr�켖��t�nUt���.���iF�h��9����c�<�$��#��qEG�u�ʔ4��0W��P����y��
H���������7��je/Pm;�;�ߠ���=/z�u��!���]�m4�7���C8���E��m����q����]�+8	a���a��1���W�B|�rY �flƻK��X��������.x���ƥ'Z,(߃�c��I ]'�=�%IlRU,�{۾�O=�y.�/�_�H��P���y{Uy\��1��Ph�"a*�l�EČ��_�ob�m�xn&��j^v�V����"���D�@D��	�ubu	(9�?�Z���b�vQ�ڻߥ�Vb���>7�p��W�
�U��V�����H���L��+�f^��F��]2�\���m8^��Q����VOp�����
��Ѱ��:cF�׀k�z��C������wax��o�3�T��@꒽�9����1~Ų
(��"��J뽡2��;
�6�-]�C)�Q�|���i�ԬX�VS5�������� �G�NaN�7�O��T|g�[��=��i�x?�TV�M�ө���@~�}��!�yىE��X���}q!�)��G5K-�=r�6G�����.��b]
�֪c�7�/>�v��!����hh�W�z>��-��ɎԬ�H~��X�+��{��D�:X��B�qӂ�'�@���(�a�S�E�^�qpɈe[1�x���2�o�L
��g��
r sK=ۢF��V�U����!�`c}D\�~�k��jү�Y}x�	��&�������Y��X���xZ�q�Tr��F��g3��u3C;+��E�t�%��C��.-�ju��!:��%��/�{�̵ u�k&�jٶd�/���u8��%��,�Sm��Se,�#��t��ebЯt�K"�+Ug�]�S�d8�棴��s`��"�nyt��r�-]*-�����x��>>R�蓯Ph ������ ���F���E�p����v�єD9g�Ɣ7:�"���Ln���/g����K��s�+g��Qaz�e[|�WY|Yzu��e�<�%�H���̿�P�50�ڼk	��I��]y����P3V~53�c!sų[��%�vЙJ��t���Vr�
�\,�#�O�8S��*x�~������w�3K(�Q���M�1����G�Ӗ�!�v�[�l96�A����2�:P(�eU�$�ZC��h��������p��>\���N臘~@ `�	\��ۑ���F�*����t߳=�"���t��cX�J�^���X��q��$CI�-c�݊��=0��Dƽd�1�$���zw>V�C��2O�v{��D"��}E�j�S��5�A�/$n*/�na�C�W���R;������DFMo��'�����������֮��ǋ~�0>U��nQO��Z�T�����
񭁓� ���?���2hMĔ+ �F�8W�V�S�+W!Gc�HM�@vc�SG�]�oF��:���M�����G��]�x��Z�����4��`k�*V/���mnq9ˬh��%bio�b#�+��5Y3���Ư�#������g����K@4w�T����H��}�Ő�䙅`ЅW�';zR �N�\���y�^{:-�5���vn�08鄽�����M4���#LV:�Ⴡ�(���U2��_mZ�Z�gkU~��5�&�E
[!]�s�.�?���x�T�p�Y�B#- �;#��ݺ��ɍ�ߚ%d�W��m��zg��r�ܧ�%��F���N�}u��M!WA�k}<8�F�q�������!r��
���BQu��]+@ې��`,D�ʘbdy���G�>�.P�_O�a?Q�[������&�hץ�g�n""8��)kM�d��c��m��0/�l����fSbQF�`�	�n�<���˙�:!�`~�G�E+o5�n�BJaK�Z���iAy� ݆�*���dF�~�=b����)�L��_�=���������oS�ɹ�1b�RT<e%��Ҋ�'�����g���:��%�3 Ƞ�Yi~�����I����l��&ƼQ�y��9U�s'�J�K\���*�UD_�G�Z����~�^�G���Ծա'�c�0ס�A��E���¼����p��8��K�WYi��;]��=$Fr��2��Kr��q����^�����M 2�!�S��+�Q�93ൂ���dz(�q�6X�� 潓�9�G:e^q���I�RҎ� �E��+������#���X��(���Y�D��2+���� ����f�*��\��C�(x�z0����[��̌��y�(�^ɚ�@1Õ7�X^oFRٻxm�ԋ ���g4F����X��A�<@6JB�{E�"8n^��G�M<���u�$���u�ZJ���9��J�,�4o�3IZS�6�	lx��*N�s����@�����G5�{J[� �.e�(�G}�W�!�_Wp�&�V`3O�6�,\�N��b ����Sr�D�������S:�n*n�U��d�k,����]	|�C�)}�~Ow&�)�=�����m�������,=0U/)0�I��t���7�9��R햝&;�s;[���Z������8�����5�h[��h��J���s۫�s�ܑMa���/k���Z/^M2��D��(���������"�i9�d���J���˳��d�"��v?����b�T�(U�J��W�˩a��CYO����A���R� vR��m���z$���bI�5�S�����V�:@�"��8�Z`Y��Q�c�+�U7�xq�.�)M�k�8�0��9ߧ���d��"��z���-1��i��C�:ǹ�����h0~�q>�%"*E��j���Z -S�~����i�hB��W�S��e;a1,�+^y�0K���9{��KM2!���{���%���D�e(����d�G��b�C�_o�\~pᜑ"m$־Mɬ2����PQ�l��4Z
�⽭n�u/5I$c��
��B��[��!0���{̉$^���;�h���])�^AK��[L��r&"����o�;�HF&?D� �����5�p37��{J�w^RȞl��N�V��RZN��9��֐$�GO�-�(��Y�	��	Ҿ��������d#כ��w��`�v5���y�$U�	<g7atJ�֚@����F���{����{�){C'K��\ƖX.~CJ 5���V��X����u-KNI�ߍ�y���wG��s�0�KBmf,,\�(r�Ü��Of�S}�~����q4���2H�,Wua�Z�
����8��7j�U�.P$�	x: Z6�F���
�I~���Ӧ��V����p��h.K�O/�]<:�ݧF~��G��S��.���,�6��ˈ�x�O�с�)�V��T�
��F�K{��z��9Pu?=/M�3�^� ���0)�hU�&�|�H	I��E"�:"�
�j��}��$�2'ijZ�7K���Fs.g4�� -t4�Q�E�*���u>�q���CI��9�ءX<+B�p��%
�%�kO��~�9�=)�L���?�Ý�[/�q1�5���R���;�w�J��g�`x��9�6��%S���I*�&�j.�A�����ѹB��%]x�	C11�>�.��c=�"�PZFG����,^�S|o6�����+��2����q�W{����)��82�Y7.��mQsh�:e�8rf��v7x���SK�?�볰�H����%�C�!e�d{��[m�Mj�#	AiV!����O�>��r��F�&����M�DJr*2����Ⲑ��s6;Zr��2zX��XS����)k�¿�i���ړ��!Q�1����ͺ��
}��9a[E\~��zda�M��^=�aJ�NL�62h���Y�5���e��
�M��Z�ߞ�o��c�	�������z+��`��><`�(!X��u�Z��j�6�h�e.`���^β�%�޵ю��������{�[�����C}!'�Db����S���s��)��ۙ���>+ba��G�6�$���l�)J�J���F�j\[����`}A��U�9��5'/l�,��.gr�wǩQ+Q{O!w�K��$����
Gq���X��ѤP��=�w;�l��S��ߙ�T��b��4�����6P��\���U~����0[Vw��S�?J5���i-��3b/��cz�����s���~�/e?>�!�C��f���->��=��7�R"�y�gy]���1�`����5r�&��3��':as��1�;�#�Y�׿�p8"~���tj���FKq�O���wL�"��vZ?GW��V��o"�P�/t���N��J��#��tB������lSw�!��;
��+ӕ��TROf�q�p�do���\�mti}��W�<'�I�&�9�B� ���zX������fS�Pd�NW�P��hw�(�ˆ{߇H*B�%�ސ6��*�#�P�J��/��!�w��|��UP�|�gcgRX-zq��E���@P�)��SL�$�S0`0���7�j��
Ć㐰%�j(���[(�I�!��J����Q��2�P��¬��Pm�������fBZ�Z��O����鸡mIi���KX!�?Q�l17ٷ�S��xȯ!䉨:a��vU�z���A%½F���;'��M�v�Q�����5y��>�K�AV��1s���>�������`5{t�aM�I��s�J��Y�p��
�[k�`4I��v��n���b���r���	��=�3�C퇦˝L~Ȗ�Ʈ&?_k���W%�U�k)�IQ��LV���S߭��� |���_y1�2����-EO���f�ų�4h�B��û�jl��˺S�c�W	�8;A/'�c��<C>�a��Ә'���WY
PA<�m\W��bG:s߬�hֲ���Am_�׺�L�WS��R;�g?}��ؿK�'�4O#xfT�:^:����˱Tx&�#�~�����0�Y�4!@��۝��}��G�ʦ��d��T� 9&��1;���'"W1�U�z��O�ތJǌ��!kB��K�������P� �?��Ѕtp[�j_R�57�j��Iш��<�Z<��vF5u�g�J��sV���n7;�.#� q�C.{;J|��a����P���y=�Z;���?}2M��K@��ܽ�n�q��y2�h�^x��	]B)'��w�*���E��߂a�~`�ڣL�M�.3r��>J�]m����Q �E�ĺ;I�u����g%Û	�,=�TS��J��w��֬��=7��_�asl�@��Q��i\;��.G� �3IKj�ͼk�)ܽ��d�IR���D��,]�Jn�&i��Ӆ��m����5�S|~��}7�%P�
��#�g��e������艁1�~��J�aM�����oP�2���j��A �T����W<*�_E=�pf_z�o�>�"on�V��ْ�	W\i=QI5�tՉCg�K@�3���/q�y�j?�NA�w �O�p���rm�2I�m@Ew����h{�'�7bϴ���}��5L�͌������Y���kG�;�i9��PZU��O�B�W�#�s�.6�H.��-�$Q��s�&��=m|���I�
��hjɈ���C���-�aEn}�?w�!��x���k��s೓�_X�7�:a�YV�c��َ-j=t�(lY'�����{�Z�D�I��D@=���
|��JP�HW�E�r����D-�q�D�~��D��?��W�Ю�*3�%2P���V�]�>��]*��tu EV0�>�D֖S��Cw�\߯�ZE��sT�ā�;̥͊I� ����og?Nq�>�'��'�K��� �2
F�����<��[OX구`K�f�˹��*E�=Q(�/��A)���tx���	���񂗃��z��8�ah��Sa��n�ֽ�Y2�k}u�%��>�ǀaQ����@ꮍ|�?_���ϓ৻jjG�����^[�ee)�u�aΒL���@�Z�g%T��YcooT~K�:�l;sa���x�1H�ͩ��S����?��W���Ӄ��ө�J<JhF>1`��B�������HF4�|1{"|������<����#�&��u��Ѯ��M����>ϵ%��B�W�C�7.$y/0�C�JK�6��UdD�o�3�]���7��.U�x����g���h�m�������j��
3�n�q���iq%��:13���!,/í%I�d�*���)��hu96
x:>��`
�OE���@o����*��T�c������,M��%���{�n|D=-�����6TTZ�;a�#�öم����O\ƫ(�
�:���J��O@�`c�ôN�IÂ� �g<�	��z���p����WM�W���t�
����.f�&�?�ա@#��r�_'*�f��I������]����|��'���TN�0��ɽ�2�:|�ر�ɔ�vƹ�1������9qT��o_m۲�tV���$����Bg�������kl���A��kyO��y�N���V3�Ƭ*�-�\����:+�7�N�1�;W=�忉�m�R^�����8}|����g�u���ߕ�;����sq��:��#,S͗2;���M�����E��4��0݅R�z~��2F�R+�V�*#>-�:%H��¦��p!�;_�^p*�1��g���6,h�@mom��2�m��ES�#�dL "�OQ5�R JT���?�(L�UF�ş�vx��W�/O���;h�h-��W��{eq)|�(���4r����*!A�kn|��sf��`QJ#��`�S�}�Icq��k��e���n�Mz�/�V�%W��G�R��k�l��M�]<����˥@�v��.�z^�sb����� /.����.�bJ�Tq�S^M!l`�A� �N�pq8?�]���*��>)jY�3ڛ�tU���K�=��ɷ��ɂ���%�	��C�p��*LvoiW�x3����h�ׄ-�� b*е�����1ǖ	mB{`��"A�mP5X���t�
3�a�g�I\EggOy��ܿyW n�#����Q8ҍ�'�m���p�O��n`/?�|��2���r������Gd!�X��+��0.������d��&�u^@�u$-�:D�)�EyS	mEI5Q=�d��7.���	W��0Dr>�G��)X����[o�iTʰ�r��$��Z�ϒ�xKi$T����F��]����T����}ܯ�\T��s�Z��YB^+���e�2�V�&�}~7�V����`���p��,���Ya��'K՘���
(z-�T��'����e��9-~ϕ���_��y�B�9]��s���ҕ-��1t->$"'�� ?���ď�]�u���GOy<��b{�)7q,B��� ��;*�m�\�(�*-��M�̄�{q�y=7$�5����CPM\�6�G���.��
jV��⫒�y�`�<%��$�)&��DkJh�ꁝ���cJ;zΠ���Zt�XT��t#?�5(�3�1AO��1�u��c�&n��GH�[�Z�U������ɍvNY�0n�z_l�h<��,�%��?�twK�oԽ�����|5�]p:�W
��@K�k�/�s樹���%'"iӍ�9��tLH�( ��?{��cf�=
d�f��l&���	�qJIG\It�����D�MW��^�<��%X���P
	mV��+�D�[�$�UT��Z��f��G�H����oBV�΋���<��,�Q�z%��~����,�>�t-$��XA�P���[)�(�G������*2�5C��t$7vp��s�E����(駢�J}��@�#˴����ϥ��)
0�9T���q���/����h�?��8�lR4���3��t���vJ�ɩk��Нz��D�H��l~�\߀�C�����үPR_��R���Jm��a�%���:�\Ã�N�]"ہr�b ?%�f1>f�� ���W�@ ZB]<.	ͪ~�	o����'-��'�6�{k��t"�C�({�7�o8�R_�/��X`��5��xlՏ9j͝��!Xl@�f��Ⱦc�O�o����dJm(��`�E�s�y�2���;�Cŕ��%�%�#m0�G,�!D���R�񒯾�F����*��6u����7�*�9Y��OT"lq�8�f�q�h
��� ����o�l�ѢU{9��J���F.��Go�����(N7�D�&]ҠR��B�3���ƇIĎ�(m��z�n��.���_b�1��!��:�]UjJ�U�V�R�m����G>NbySs�U��� ju�P?@�\���+Eum�NtC�^.B���IIQs��#�Q��. �iq�5�"�[��3����x�b�I,`�MK�Y�]r�$x�ӡ�|2�҇zp�7�g�
�ҋS���_s� oo���PJ��E5�bW*#�ğ�Z1`u�$����u�����u���/��>���v�-ǽ�W�B��y�:/���cS��#!pm-)�лҮ˷%DNd.���x��8�v,q9�&�^���ÔƫǍ��X}ӻ�8'?z�p���V���B�60���������{��:/tM��+=��!��˧��	B|�,�ofJL�x9������1O�`�`�'K,m�d�'����fk�fGC�������L���J�at�߃%�U�ڿ$�f�L��"��{A�����t�}�x�'��s�RU^a�N��B]��U�q�:��:����'����SJ^�&���:�ٌ�_I"W{��P�P�q��
m$��@*���A�q��6~����p愎m��!��w���Q[�B�3l�{ē��0�w�.pc,�j6���"�`���l�M�ﮋ�9Q@
�7���)�ϩ���!�=�`���k��5��Yd�N�lb��=�QU�3(�
��g�UC:�#*,[w�q�ɶŕ�ܖ�8��#�$�4	��8J����'��J6^sGU����VH�j��"I��B���Ua����M��0�����H���x��v�B ��C���D���������Q�2"*��;	�TE���HM�s�
�|,z}�k��8��h����v�ZH��m�2��#y�M����G8�3&r������0��cf衬��|������O�r��[�cpHM0�;�Fb+C��㱷B��/BG�QyɈ�^����Śg�|�6�n�cM��lg�S��ڷ�Q����n��ac]����u+D5���5�*��`����zu��"x�W�ip#�$l24���0��T��mM��J5�a�ep��Z*_cߐ��|P���K���ȣ�ֹK;��!A�')4�'�dR�űՓ�sV��벾5)�57~EgRd�
-ē]��(W�ȁ�YO (d�W��3��\�4V�C�{�*r�1��F2�C��1��}$�P�]ۧR�5�M�&�r�X�QM���L���>��X?k2UM��
�Ba�[�Z�O$n��kѩ�5ګKLԫ��KM��P��j�vK�>Q��6���\�C����w���օu��;���p��s�1胗�T�ey[�H�M���h|F�z�x��F�0�G�0Cup���3^���y7E��Z�wI�M�aBk����[�Wԟ�\�ݶ�3V�"�`����5)^�lW�Q&�M�E���< �����G	Y�f�%6�R���?ˣ4�x̕#f[�J�2Ɓ��Qyؗ���]?3Q���--��3�|s�)1��0�k��8V$��
	�	�o �p��_�{%����cn�r
K�i.���N,i~rv�����v?�r�YlLP�߹�]��n�*�ct��B��Q�6�9 $S�H�,4������5,�1T|Mw�BU>��53������z�ۻ�y1��C�����`�`
}ӽ�V �x�H�~�t�>��y�e��IUdͥ�a�~�R��Y���?�'�Ќ�Ԋg�J���#�����'d?����n8?��f^����$U&����H�W�+h�H�s��r ^��ϯ
��� �M-������v
e5�o x�=ǡE�E�Or�	�0;W��H~�3l^��(���Ԩ�JF����u �Y��s��L���@���L�.��"Aly�(f_�>Ro����3sf�;�s%�:�6i�n�ƭ�y	������� ��c(�E�e�ƙ2,$�bB�!#�;�[Q�-����=�]�g��K�U~�8(Q郹aD?���Nˑ���ې
+�f���g�\"������������ȟ��B!�I;ޫ�?ƍD���x�������h�������=֚̃�"�f ���@�����������ˣdur�n�n�RIw���0봊. Y�h��A���~�FC��|���b��:^,t.���ހ���������
7`G�2$A3��?Iy%a<*gõ3�l�-�`�!�ʹ�0��#��z�hHOW��|@���M�pI#�E�n�u�?~.b�	Q����~�����ߘ��0��.�@J��2fC����t%�egAW�����L8K��a�ue�0�Mu����c����:���Y�2L����9(u��:8o%�4�[�� �@��r2(��T;H��PU��|�)�%}�F%�|��3�����"Wr�_���Ӵ�ZFkH���� �ڍ&}'�p����a���>�J͍�G"�!~;�֖B�ah���s��5����s��B�x<���<�]#,�=U�w@%�M��򗐓?���`"���烬 ���8��Fݳ=C�Zd�@��q�ʃ,{��O��8�U1a��W�'�)�k�NV�9�d�]<Iu��V�8����R�+������ԗ�x�:�'"4P�=nw��L�$�h�>M�q�1�|�A�wz!R�R_�iRߔܻԟ1Ö�q�0���s-4�J���ڿB
*7��L%lޯ�OR�`�e�c%K�]Nq�̛���:���ԣR�G{z��L-s }l.Ķ4q'��)�a	(�Ă�$����	�S)��ަOgc���Jq���Ql}�S�:�C��Vtsv��f�c�k���,��J�zD��-��|&[��:2�ɷ�m2��rMc>�|X�Mh2��5�A����4��*s�>�8�΅*�=E��W�=�{�s��q�@ƉC�kX�����o�,[��G�B�4@_���#��q��V�[\�N����	���˩���F�!̗���r�M(D��!>f�8�yjGׇL��D�
���mI����|�	b G+�/g��a[K����-/)��.�����^��!�M�'w'(��Qpw��cy^z`|�Ȃn�j"��܆eRK�:�Ȭ��Ͳ�t
�5�1�16���L�����,�~��β;n��1�J�+���'�_�d0Zx��D��� 8Ј���^�����N�#Sg�8v@��L72� ��l�f���v�M��wOm�f��:��}���gI�ż�ͽ�׷=1�.��=��1:�ymb ��+��#Ń8�'~�%5Ծ~��C��f��:�&V���Jbw{"

���g�[^$\۷��}��{�1g�=v�iTl���D:U�G��dec� d�z�ϙ�M��d�H(�
�\�u�� R�$u�6i	��"!U0���j&�/��f7Whz �}L�3�8g��-Q�E��IU����,$+v!c+Ȭ9�����N����^G�]u���4my3������/�.����o�>�>s��Z�������[�-W��x�S;�<���A� �F�5:A�J�/N�O�+��ɻMWQ^���+U���F�Z�2�[�m#4�o����®AӗV��=�1O�<]D��~�����>��0�3~}�+L����/ꢽ����I�TlO���XĚ\�[ڜ��h�A=�����>�%3���x�$��a�&l>�iVl.!��%Ը���o	����]�d�L��B*إB�b��`up�Kh�Ɍ��Df�_o�� �A���Բ�Ai�M�,X*�����+��u�v�������
����0KD��j�9vC�<��2	kY����|v:��d�3W�ցꏙM�z��q*��=�qs��76��=�[@��-JR��{y�F��R5�c���F�kSp�"�:&���L'�W�H�챲E�4�	0sv���r��$�^�awSc>^�Oڗ{��ڃr�ᗩY3�AH#R�SBqF����X�cZ�d"�=ź6���xj�>�>4bSD��>wB5x�PI+H�ho�_�65=��������)�3X/k��gQw�s�}��������f��<��)��7넷"��MW��tWh�@&��2"��cÃ�6Fto��!�w8s��]Q����[6��,:����E�kTM���k@���GPH�f�&�([`�=�*�N+Z���4���9��nEYgȒ�P�u�q���	�<;3�Fz��<i:�Z���I\�&}�qg��}C���ݚ.�q@5�����<.Eږ��
;���T�r�w{���naLf�t�(�T�j^��BB�n�LH+�*���i�&�{�. yl#�4_-W�zЕ�������݆o`Ő\@j���Or�z�ҟU,7���w����~�w���7���d̈�h�o^ޜ1��FC��	�+�?UKw�����?�a�D���F����FV˝��U#��C�����\nz��2��40��=d+*��M���@�c��ɇZ�3�詪�"����Z�gT}�q?���G��^T�H�����;�p�m�u[u�3ۉ�m~���8"!��|��I�m�RB��Nw�&2FqGjGYs�6ӵ!	*.��q�}Iʋ��5X\޿�M>�/��б���K�1��3]xIoX��n���>Y���_���{�m�SΪ[�_�ϪeL�I��q)<N~SA����j5���(X����fsbz�NX��mH�o��R�j4��-��P?h�YW���G��5U<&�X�)[\�j��>y�k��d�,���~7���#����~>pj��:�aduJ�*醏�z��,o��s�&g����N��N�N2�ZVnCx����߸����,�C��5��a��c|�u�\�736+?��s�����!�f%�$�dƅP1-J��Vxi���L��Ԋ��%�zE[a�X�L��)}���a�ն�(e�=u)�\���4�14�-�BW���� z�������y�(I��hh7{��h����v�����[���nl�|e�r �H��7�_��1O�#Xc�dL5�M��Њ�#����4��Ĭzw `��n�\��3ah[AHM���!z�k_��0=T�G3�->���^���yt����%�����Zy@>U�������n��y\"KL�$ܮ~��UG
�����5�4ID�n�t��Iw�� �Y�M�ax���5�פC�{��8�1+4�\U��D�M��-����{�T��I����"��s�	�9n���t�K>�=���L��[���n��Y�4�/�V�����F�]= �"�}�o��5/ύ)�Q'LDbMw�/#4��Ya�3-\��vw5����K��E�g2�8V�/qO�
Q�g�D�s����Ԫ�R'���cT@_����������ZF]����H��hҗ<-�ʗ��C�;Bsn��Wy~���\�k�x	'{YC����@��YjğC���F������9��)p[a0\��_��VB��(�ЈQ��<o�vFuk�i��Q���Iʨ��\�_҃��4����ßl��h�oD�*�!����َ��&=C!�ڶ��Υ�XU5�ˏUan'm�`������JK }�2���c@�Ԝ�^�E2��+�9����J�֎}0���j������/2��g�;{���9 �1'��!�	�i����bPqĕb�C�xul�����k�J����N�E�^u�8�MM"�o�^��?�u�%���{HR�)�'�h6i��/���r?���}�#Ɣj��bφ/�n���\z)ֵ��0�������f��Yx�����	j(JTP �����y���:�A#�\`��
�$�wb�O������_��O퉹�^.5g�D���Hh�u��hΑ��L��y���)���=��@y�깠�t���{熩�Z�/,��Cq�cJ�������?i�w)���*>�����{������kQjV9�uȏ���͵~/j�5mT�?O��ѨXM/�ɵ�J`ǝ<�1�q`߳����f�ZMj>�U!�u�\�a���%�OF���c�G�� �(����+���#�s Ux|�9�I
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���۳AW����{�u�)̥�d�pM�y7�w�1���'�"��+m����Ԇ�@?D.�#���A��ey^�??fi08H�w�%4|s�.���`cZ��wʸ�0�h!#k�a,�ˑ�lx���\�:f�S�W��n6��|�Z� ���h�i����fJj�Hɉh�7>���Fwyg���	��CfZCGt)�r��Z��j5Q0֨F}읁�eU9nٔ�D�z�����|sn�;f+�}{z�H昻@�������r)6�ej,�	�b<\�_k���5ȴ#�
ًr�����{�����LU��r����r���).�L���|9P��-����yet�/�=3��:ѤR޵��y�lb������7|��d�r�~�P6���c��bs�1:d��C�D��SE�_�m�$�����Q��ܡ�wu�7+���eT���˄�#���8��n�f�xu�b&E,�_�P7��oq������;�}�V�	D�
�V}f��Dp媭ڮ��k�C���BaJcG�M�)^���XR�)�,lwM���`/�V�q�"1ɀ�� c�aK�,ɳ�X$��X�r;>��5��K�}�S}�/�y��'v�To�M����Ĭ�)�<��9E\]�nQ��/f�*�
(kWS���6[6̀?���-$�q�;�Xt�?��{!�7g.����17�t���d��&]����"ɽ�u�<��e^<�>�r�L�"㐦��g��U2X� ֘�/�oD?�����,�K�����M�t�@�\h+���뵆x����k�w6�Ԭ��Ċѻ�WQ9��7d:���zN?*�C����:8$>�Q����Zm��`�A7Ɵ�zDk�C�����%����kt��-'� #�t-4!�J0!ӗ�8܂tk�;e6ZT�a�Ѝ��&f�]Z��G6:XY%�Nִ�i2�y��B%ݼ�ʂ�o��=h%r�}�����:9�L	Q ;�v� �K�ր[���M����"����.[v�͙s�xX�����f��U�S�u�3�VҠt-����^�B��u@$�e���I�r�/x����<XJ��K�Ўп��f
�hց��rw�
IA�t,�����8+2Z�~-'�['n�[bt��f�Bg.�+:�lp�lz~����FL %��l�5�M����O9-5�f�S-����[���;�5���̝�Q��}}���O���,�2z�:�<Jc�p�1�O�W���!Ҿ�X@���45��HmC/^�3l������bD��$���&�EF�F)���բS�09B.�|I�Qo=�rM�_b7
��v���Ac�T�S����u��^��AۉP�aE4}7��!�FP�3�`�M�m^��<�\"��Vu�E��>	���`[����Տ1S0cx{���~�5o����Z�@�A�[Fb�V�e�L�3㸟�z�mr��Mȥ�$��XV�;�7�D{A��� tZ_�>6�̯7n��/���.ҳ�I������;L��%��`{c맖��H(��.$eP����+���HB��J:�ި!�#8�)Nw�vT�e��H3���0���~dJj���ۤF�0�/���XػM(�M����{Y���5�8$�1MOU�O��9�� 8ל��	q{Vs�w�|�"y��
�����}٭a#*��k�?.|�a��Ws�xoj"M!�q8m�>Ȉ;�G ��q���&8�5�;�0D<r(���I˨��s�r�(z؀�� ��4��zZ*�
�X�֠Pn����ۛ����j6�~�z�����?ɛ�����@> |������i獆��[6�Z�P����U6������Ξ=��rK��,M�:�\�� *S�*\;� dbz>�gOl�smn$_�o�	���/���%������R�D����R��Xgi����o[��P>5��t]�.�O�������zNK�֊�ڍ��%KG��|?t�E<�N��{j�����V[�pcR��8��͌e���TM)
�+����be<3���(�k~> m�e�GM�Q� �h�V���U��H�Z�>h��(O�uP�i�%����c�־��r�S�>&�7����-���צ<���5j�AŪ��7��y>_W#���2�M�k����;��XVb� B�����6�x�տ�6Q�NM�v�Ovn����6�i<oN��Eɋ���v&Y�v	���~c2X�p�&I|y~&J�C���Pd�n�i�d2+��8��,���ts�*�{t)�.��w�/7� ?g>�����z�"m�`��{f�o)��Ϸ�����١F��%?�o;o��&m�)�[��2N�O�[����[��0���,NHk��]o*�����,؍r�.B�(�E��
��6�:�Q��k� �SE��|�wP���ys5?Q>ա_�D�l��bYj���S9W��n��ɖ�2�����o���o���D��^>x���c]e�Wu_T$9ʁ�_I��&<U/��3ڡ���Z��jq�.�I�7���ah�a�F��c���i�!}ie10#�4c�@
F7���!sF��PE1:�ѿa-�q�h�E97y�n{���ep㌊�E�n���ʉ�E���f(:�e7�[0ǘ|x>^JF�� a�ȸRؕ"�P��"u�u�M�������7�q�LϸKϫy�ui���y�!�O����P�o�����O��SW�Z�Ss7_��Ȳ�7p
T�ֿ��>������r}���%D�ߵ -���!��ű���\ƺ2wÔT|K�̼�64#�t���@ZQ�'	j��Ұ���v	�;��D�׿J�٘��[���:H�bg*��`N!"�ɲ��~��`��X��$�f���*���J7��MЦ(�:�U�O��H)��}��L�뉵��2�s�)��z7��؎��V�+��Q렬DrMży3�^!�vF�a[�~n�����A4�-G%�7dT�3?�MŢs&��Љkm��m��y����?n�f���R��_��;�QK'J������#6X	��}L�y���c�L9��ւ��`ۦe�
W?("7�W>>�i?�h�-�Z������
7�2�I",�k���h�fȼ����>�tvf�KM��굂�T�sSʾ���9|N�a����=���cOk���K�C�r��t��KAO�0>r���t��`3�.{���W��G*̊��_dg�+Z$�)�D
ʡJ_L������{��V��K:+S�����
�.�1��O��y��	�j{�F�xӸ�}�H4�|����=�?w��o�,$uݵ\T���Ԝ.���t��0�h�is _�TD�����H�l���#L�f>������H@-�̈�_�uH0 C]���8Xr$��m*�2`�y�0!�8�7:'�q'�0�K�/�^IN[7>����3�(�jw8�*�I<my q#���H�.�e=`��ǃ�Ui{��B�߹| �5%HX�[-f�Z�H^AG��(N����k⽰}6���9��K<3�������<�7��Y#�Nܣ,`F���� ?h������Y�4���k���!ADƖA��٦�m�7�_jbn��h�-hN}�gޯ"�R\;I����XCI2��܎�,V��MuT�P���֤��24�z��qR��Fik߉������������.��3'ג���:�(n�ћ:Z8㴉0`J��ܝ���h���g�Y��r�� �cztEU+Ǖ�¥�FxA/�$IPY�v)����Ud��v0�{;��3�ز3	��үz�@|��ag���_!B��t�v]�vU)T����i� �[��{M{�cJ����1�H�U�h�����}���e���t�G����^/�����J<=��z��l��L�H�!!Ι���4�M[�Y��|���cp&#�U�K�m\���/��F�@�`0Y#.�&\"����3�sSv�{�P�LY�"��fF���%Wq����n�`7<䷣�&��lG��B�rZZ���\
�&�О>)�iٹ'6U�ˑ�:�BB��F����W�8�Ȭ��>1��#x�'W}{B���;ߛ�A}t�X��f�/jh��?�PS�4v>PRiJLy	V�d�к�cv֧�&�D�|������f����^ U�)I�9�V�Ǚ�u��(�L�h�
;Lᯑ�Eu��ؗ���`W#N���L���X�6�]��G���w/�-�%s�I�2�1�zi��7�FpV�PP�y���J���.�,4B#��K�:�r�Og�ol,��ڲW��2���o��f����=�Έ)�S��&�	��
����<�zs.���q�VF�`��~(��)���bB:�-���(���c4*+z~�6Z�--j�&gR� �3]\����م^'Vibz>�.:�B���A8��|���K�G��b�Y���;wA��J�^���*�8�� J6�1( ���;�q@T@0ս���>υ��l�RGxz|��>�஌Aݯw�������q;G!��&v�͸����	l(�L"�LĒ�~,/��Z�f~`��[0��.��D=p�.=>���#k�~�Xh�]�d-6M�-쿚A��K[�/a&DTl�%~�=���ݧM���o�oO�T;&�73Rf�;t|�L�ԙ/ڬ� ���u���c �*�����4�n���s��ɬ^��܎7��<��m�C��25"���D-���x_�[��x����-Dk-�k�$�e�hx�A��Azvy��Q�����j��4.��yz�]CąB�b�~v�<��9�7�=��>�Uδs ��v�R�S7o��渾��u�m&�$�����@��䈛�U"�RyP���+�e�����)�Iw��wPו5�i�q|���Ju�m������m)���#a�)���-�v���Aq�Z�c����KnGΩ[l,�?�U�u&$�t����h�긊��k��	��O���w�%������g3�yr�������R���@U'�'ΓT�º>4��T)r u�Q!qz�����]��>�ZM���˷d�O؝�n�BB���X�BL� 釞Vqf�6Y���;���L���u��)&���hĔP#��	އ��\}r�3V��x��"n�|��M�� Fb[x�������ll��¤�#~�s��q=6�L|қ=�z���[^�uo��+�p����h�����J�@�r�oe��Qc�pc��Nŷ�`{�ʂ�M��P��\?�w�=l`^ӧ�HM������&`��,�=w\��q�H�����Ư�E�5�Y�0��Y0�;`��ܾ�
��h�c��*��u6�H�bs��;p�ށ���n�=�:�D��ڵb�S���?����2�TZ�&�X������ʛp1�$�$B(�8>�i/��P��*�#g�i�nx���f8� ��A�n�i ��A}�[=��z����iV�I���@(��9uD�q�?���с���%���ˍ�J�Ov-ơ�{LTV� ��ePn���s08����A��{���ڳD}�%z�߆M+�W҃�Gp�m0d/�5���g���1���i"��F�]�. wJ�p�A����v�������8�����'�rK_/�퟈����k@�}��6^�@��f�N;�ڜ�J���	���1�oc��`҇ΛP����	�F����~Oyi"�������ͺ�H/B��6���y��헠�C��FH��;��� o��nUM��{�6yB��zb.7~�m=;Հ1k����.��6T����8�gj]m�e�n�'�AI�d�hh��0<x�Gl2���İ��}|P;�������-B�`�hS�X�M�v�,lJ�t��E�Ťu'V���x��c�y������g�7�� �6�i�}{�b�3PU_c�&��*�_��S6���Z����'
��Qjó�>�W��ڷY�O�wRa��^c�����B�����p�deѱ�[\���7�95�x�Q�E���&�H0��8�1,�)�㯍lw�M
��S�l��e;(~�$�K�-G;�JxP����"�m�u}sb	�l��{�-%/��tj�O�?�!m0^��)��y#on�K�Tr�٣�=*����Y�h�e/�D��m�E�`����N�@��Xӊ���?@�h��q�"�r�����李/^��|5��L���a{�:������rmc��(�&Q�<�'�k݄݋Jeߐ,���ʯX2���� �O�G�f �ً�-ğ:Z��槞��c}�I#.�=Zp�}��G�~��5b��-�_x�5�%��f��*�#��ή4��L�Ҏ��ڤ٭�����mu�K����d���9���C_����T�Tªp�8�
�>rz���2�o�b��J�h5&W5��3�6J֓�7�'������O�	�_�%����D�C
����#�]�$h��,u6z&&GJ��ɱ�f���!�Q��ۛ��A��2>�%�VP[�s��|���1����7 ��!��^<0�_��e�?P���f���Hg�J9h�8�Hb�q�ɚ��/�R����B��/v1<�:"�>.]~���.`K<�c.�U	��T~#�Լ-��w���Ӌ�n`,�^0Ӧ�s�D�>�M�����@`Ҵu��/p�����a�$R3u��b6表y��{0�����ז��F�E=ַ�U�H���Xє�X�3��-!$����s�hL�-�&;�@Cߝ;خ)��z������F˯mt��U��He"����uY�=�dRK�S���}C�}p�=�pę��7[��``d�PT�ދڎ�+�a�k��_G_�i:H�V���f�Q���Y�}����nN����ޑ[X��"U��ob���k�kSݵg͐ ]����g�
i��.�y�����Y�s�p�㟬B��!7��"�*�����Z#kӿnN��m�
R��L����4=�-)Ϲ�>o���j��7V���-�B�V��}�3D%25����+`�cU��h#$��h�.��5��G��Y����`�d�gd��N�H!��>��έ�E�a6r��T�g����ka��Y�Hge9V����T����5�k�@nhfH`�,��p$,o���P�O'`�ܖob<i6��-c�|
�m�cg�񋈣�'Y?_U�Ndh�r�vkt~���Q8�7�$��,�#3�/� V��1�N1�5j��
f�C�`��po:f@��X�Y�[;G��d������B���W0�b1C�p�d�W\�I�%�}�z�t�ܝՏ9���<m�N������e�'�9 ��7Gy
�./�dA;���"��2��s�3X�[9Qu������dj������S '����([�� i�4�
D�,rd�p�EQ�wZ��o-U9��P�}����	ک#?�Q�T�u�GU�ajI�>2n��g�cO[@���q��o��Y������tN��}$�c
�3���'�Y�;zM� |�=�NI>�@�1HUx��Jsa`葲��qPd�S�;�9�C�y�=l8I�+���ٴ���6�J:�X���'�b�%̪!(�f�Ě-�e-)�ՙV��B��6���<��^�m"�w��f��������D�� ^���lc��h�7*<X� ��I"�p����E�J�ʷi��ic��yQ��hH
9�#��{N�I�@�m�#����Q�~,��4]蓖�5IE�+o�q%�ۙ]��s'5�T2�q<Yh�0���E�Ý�M\9��-� �7�S�X�7�1�6��/���-yn@Һ��?w�i!�Y���ത�*Zl�E}��T̝r3n��$��)`F���+T��HѺ�7	Y3!s��kZ�Ix
O��Dw#������"v:��ջc-e��73T2W2SU���^t�^b5�����,� �~�8�!ײ�c@A�a�����m����!Y︨���t9�=�@�"��9TE��e��/�;�ټ��a��̛�?U��r�{��;?v5=��R�C$*�0���$��"�G%�9y�2�9h� ��n�Z���=P�r�Ps$F���G<�`�Q�@*�M"��R�D����	~��I��B _���$q��E�����%��M�XAg�rs6şI����=��/IV��}��VF�:z��-D]c��:�F�zj]�0�@Z;�?����K���$�D�\y��{�B�d�~��z]Dpz/tH<#.� M��C���V�Gg�
<����٤���[��*�e�y(�ǡr�qo���s�#�c>eG�ze~���L�&��]2Y�4ى��WI�-��Q����B�>�+t��:VG�γ��.����;0uo!駬/&�����o��J�w-"O�� ���c�F�@<�'�ݯJ?Q2xI�Bx����X�Z��Ӓ
~ w
�0�	ݠ�wJ��l ��uF�z��r!��-=�Zs��G��g���Bk �H��^��|�uTB�k���������Y�K�g��ůranο���`��e�@��RC�ʢ�\��{�޹�Qw���EP54H��0SF3�p��kaxcӧ����ވ��|+����e���ŀ���W��m�����̣��s#���R��nu���_}�<�g�P� t���x��A��[�e��5)2
ZQX��P���'��`+N��[{�p�J^��+�R�|G��Xp���������
��l�N��
�h��k����W��Y7$}���
�?;|��ݭFh)хٺ�Q����R����h�7-g�B&��y�'"'����~�?�71hOF;>��r�	q�6 P"sTw���gS_�Mx�����"-C�_�K��j*L�L��zRq��A����A��P�x<�u�^��''�4j9I���$ݾA�@�m�6�m���Ҁ��-�M��?�sEG�ē�b��t��#�V{I__q\F����{;�4�aZ�@R�����/JJ!M�n˂d���$�mr���5�ٚ5���u�x��T�i�Ynk�J�cR�։��9�}Fܭ�k������"~bE�ژ��x0��̺���`#�Q�����8����Rm�+�x��yܐ��<w�q�{�nz���[f�+��C���g��������O�?�O����]����r�>( ����R�g�o�P���࣠����pΒ$��-�mO�U���#6~�:}�qߓ3�<t��P���X$�����#���;�;7�H�hM� ��������Mds+��T�����n=�{@^�vL�ݡ�'�`l�Ԅ��-�X*Φ>���?�gr]������*���\�4?z}��L�l����d�M������P��>��%p*ULߙ/��H�?��~}VH<
�3�FfG)���d��tԵtǵyMn�B�JX�m��} �ٓ��q'��f(V�:;E�()�e�ڟgIo)� ^2H0Y0\w�\hG���B�&�ͭi
�������,(���`����.��Th�[���QFb֧}�P5g�Gh�s�u��j���T�O�b��TjS3�+�*C���i�'�O�+MREFծ䍭�$�Qs�zFf�6[�u7��n��e��JC`-N�	p���0��82�|67�:Z�i��.<{}��M1�a�n�@���^;��$�q���1^fxm*��6]ך�z蚙(,Z$���EN��\1��˷�h��<��f���I�Fd���p�&�J�����2�pK�W;�MJ�61�����]ܨy@׹�c��mQk�����2|9�L#!j��x��$�����8VM�����LN*Z�3�]��X����.&��u{����&"v������V�| ��9.�J�~>0cO�����#�+J]�epB��e}Fq�]膾%��P�N���hbKV5�U�u�T��O�s��BJ#��ZV�TلU�.���E�$yW3_b,�=`����zYAD�=� 2�[��(ݎ3�#�
��ªQ���xJ��3j����fF$?W���'�"�c�E�x-B�@d=�^��2�sמ�pO�:��T!����QɗME���=�A?F�Y�	h�_�%r�@A��ߣ�A�-�c;�@Q^ӭ����X��y���u��M�mW���vIs���d���5�;��d��H�����h'L41���?S�����B> >������?�m-�V�;�Gv��y�'����y����7��o� XMئQ.>�2��L�r��.� K�C�wW��ǥ*c��A�Bi�6+r���!��I��v��j���� �n�.ϱ�4`�M�T��أ=�O@��V��"Lg�T�m��)/8���)zL�����@�K1�i:��]�f<�h$��
�Ք�� ��nv,�R���� d���\�o~� P��D��-����
�S]��KY��w�h�������$�{ޤ�����q[9A�z�^��ŷ�3�n0c���ϔ������j3��f⩪x��j�x��5r�TN4�-�.��Ah��1�[�p��9*�6��
���T8!c���4?�Yo�aA�l����þeO���<)S
���@lX�I�1uGF���9\��~$ ���@�|����:��l��0�Cv��[���iR��6i"�pN޿��0a��'�4/�{x/�1�� N-"���X7�q̊���j]��5���)��|�H��\|:�n�����K@�Ȭ�`5�56�9�0�u����[+�I�e��37�"23n���?D�LaY��Z@#]%'%�B-�9h"ķ_��W��x�H�k��Æݝ��K*]q$P��Y�G���)�})���
�� W`9󸂈^@.�5��`������S5���j��A�W�f�W�l��SD�l�xW�P��)�x���&~�:u&�i�,� fs6�[X�a?5 ^���vF��Q ;� �.�D��3�lШ�	G�������8���v�,F���_�:�3eeZ�s!x2��o�P���[�9Q3�kŞo�/c�9����ܬ�C�!�GGN�Sȹ,P`E׮&
����\/�ŀH5㡶bL��8!?�Ή^����T:J�{!H1����;�IԦP��oJȷhX�r��ڰ�v�n)Z�� ��zk@a%�(A��g:(�lqEܛ[��&��73�c��)�,�\W�#]SZ3���|>uK���	�*�d;�or���j�t�D֛t�7�j@ؿ���d`�2�]�3��ع��L}�L���K��Y"��N�޷���_�����÷k�\rB�lU\�8Q0w$�ٕ�	~��� ~��❧�A��@ap� J��������o��=����Ve�n�l���m��w}�_�h=�T#@i����Wf���Xl�Bs���R��/|���0�ī�zO7��$�}�x5�z�ө�SCP�61�u�rxuy5�t�G�K���$�D�X���N�p�[����+ �����Q�����~o�<����w8��/��ht4�pL���jl2�l3��Pi)��Յj�j=IWr�D��8x�fuȮ"R;cB�Oh���:}\1�H��R�3PC��v9�z�G/�����j����խ��
�)��:X�?�k�`&U��o��F��>�9\}U�Д|U?�����@�*����^a�T7+�H�l�H���'w�tۿ�752��Vk���v��,�6�H����m�M�g�|mϳ���fjP�U0y�5�H��n�\S��Pޝ3���G��Ri�V�L����W+��P�X~ n2N㴥�����L�)#ffs��+j/vH��eV�����w��ҟ�����k\b�@m���#.C��!��PCL?L�ZS5� ��`��Y�a
̂@)�n�й� _�N���2�(�I��p�u�_F����Ss(�8�K����(ܜ�&NEɷ��W���5����
��I�N��(�Z1�ݏ鞙1٤ �OV�����V��[��=��*�A�cx�x�K=�µ�
.bm�&B�a��ͭ�ҝR�V?#f$�4���_�>�@�W��75A,?����c��!jX$љ��td�uާ*�a-���R!'�>�eU�k8�r\T�$�T.��&��r�-qKm Co>x�|~�<�������| ��L>Ӓ^LWL�V��W�2���W�h�t�cNtn������x��6�qrp��FШ�7y�'�q�q�㉥��(�bY;�9��n�2՞J���dj���&��*Y�(c�x�k����B���=�h�z�"x������{�����,
���,^�:���ݯe�Zn�a$p���� 	��������JyGƯ����C�������.m����ˣyM��5�V� {c����}�Uc�� /}�C.���	yfw�m�� DVA�����hGfL���L;
>な�ߡ��b]B�5�G.o�:��;JpE��W*�l5��D��oǥ�\���a�nS�ӳ5�����*u���{�
��Mե��S�Aeў4+��li�����υhtT?O/U�T�h�7�e�r?��Cb��}�;F�W����$���'��� fՁ����؂1nꍐ�^�����[aG���뵋n�j���n7�l�[:4H�@�2h�1�D5���y�/f�ds�8��؅�i-m�_���n�f�nM�2DHh݃H�AX�Cb���9P�[Jzͪ�ތ��x�IwQ9\�Ɯ��}2������0�V���� Jr4�ӽ��/�#ZL�w�#?xO���JdA+�i\�HE���X-<�������e���Y������� ؇|CfS�#f��q�I�9Ɋ�2�����䖚��e��pi�X2^�3R���h]Z�ɾYK��8����ST���n��$B~�җ1��~���X�w��@C��h;E9������?��"�%�jJ���>8ǜk	�3�4>��B�q׎�*v�k^V/��sý|��(��F�6�(��	1���ʱn�hI,�3@�+C����Qg�S�r�SH��iܣW�͈�!*\=�A�V��@%��؛rh#qb�V������NCCC6��ok�I��0��}=�ˈ�r��a����hr�����n-�` pR�/g���-�������*O"}��>��J�"E$�ǈ=���'��Jy��JR� =��t��!�~��l$,��CLڴ�'S�{j�	�!V������6aj�IF����q;a<8�j��p~����X�N����UA�T0?���Pr-w�����}"S����Lv����s��
���ls���ȃ�	��g,I�F7��F����������8/�c�S�*�\�3zW�����|��N��z+�	ƗP-Uf\�w�A�v�E�E 4�������3=�x2oд�����\ĩ���
,�[2�Ʊ#ǎW\����%VM�z9����K����I\L���g�#�D _{�Bآ�ƣ\(��)��� b��(�e�7"�G��Pw�A�[�����,�#?CԼ�W׎G!��^�"�A3{�CHX�H����J�� ��@1��� p�b�8�c�4{�C�u`�r��� l��ʧG�@h����daC3�Ta�&i(�xIK�1�~��pQ�CC:�tt�>刿�h�U�4�4�B/�P�����k�qe׌hR!��g��}7$�"����9db��xSa:��>]x��A����hZ��Z!:��j�E�}�a3��1n�%�R��$5�3+��s��ܩRϹ��	[o�Ni�k�tI7��@�~eYPӉȡu�Uº�G6��0�pcg�������C�����Z������)V�?H4�qٰ�l�2�~������,)d�f��� h����v�8}Օ�o9"�ٗ�Xe�/��C��GUny�'"��d{�N~I���j=Wҙ�����ѯ���.z���T@_']�i썣��<�	|g��YEĂs�8�OBX3#�EU{}�%��?��Q����xdd�eJ�l�����	���\c��K�o���;v�Z�͘��9Z֪�r�L��*����[�U+,|�ËjCS�*� =�]�O��lkr�I�d�?k��c@�J]����n��*�F$e�N�&؞�f�R�G� �ʽ �c�g���x�q@�ͽ^T��/��� K�/������~�o�X���Ah�tM��y�F�wŪ�L��UXO�r{X���(Hw�r�h8�G:ۿb�RX(�u�<��U}�@�D��h+*��4�C��ޛ�{k��4q���.ȋ����f� �1K�X�!S�޳����� ��mB��ڱL�8:]����K�P���H���k��3/�s�[1�Mng�����~�^Yc�m@HS>��r���>Z�P�w��E?�<�$Q�l�F��J=d��Ǭj�q��`=}��uT��ci�ГC�8��#8�����b0IJ����%����?��3&��a?�xt�J���]�~ w��
A8'��j' M;��3�����P\S1��0��ho�p��UkYX_���M=��)WJБ �3�jq.Y��D�DeO��PPH�I|w����N�Ͷ{.lvFI��EqP� v��9��`�)�'��-P-i*̩�e�-~��}
��GM�ynUVN0�gx]]f���"V��֖�\yZ؀���7�pgZu���P�\��V�����M�i�r�����f@c�7d���tr�%�5)`\�V����~�WA���A�In�Q�L��<����MT[ˮ(�<���L�!<Ā�sX��QjIؓ�z`�-Ečዉ�~�,��R�I���_<0��^bob����8W2'��IP/��X���I�PȒjf�������'��������b���%~"�TN�3`�U�]�wi� ��bh!��z��'�rܔ�U�Zg+B�^���m�I���$ȳ�P��i��4�N�wq%�5�-o�����񊊤?Oy�\O�����2[�z)�VuX��c�
B9㶐��B2�?l�t���O'vz&t�Ԥ�`$V�UDI��^�Я��nf�_�p�rwq�,���M#�=���L�T���	c�Α�7���h�����3.r�2�28���9�k�4(,s(
ƨM=�sޒ��ٔ����� �}%reZ�Q :��a�+>��Ġ����w��kV�b|�
nw�F�]m,rdVF�io��l,�x��Dû4 .�5]c�Hm�}p)k�w�^��¨�k'|M�vБ���EG(��7�s;�V0�A�H�X� �Su���	��I��M��">f#�M��>���b�7ۇa��!�L�C�r��"8!�׋���yk�s�רv���)a��Ln#��2��:�IG! ��qkN��⏃��a,��E�i��g�>��PX�%ϖ�q��(
9#j�i]���C��~�Y�ڧ�5R��WTg#�߄�6��pi�|�<w���c^�D��)�3\(��C3�����	;T����Uj�΀�HC� -,��Gp�⫩��Oo���@�7e�p��ռD&����~
5$�������b��e�Xvk�z�f�[��t0'$�U��9���
���5���|ܢ��ݐy>�b� ��~���0"��F'�!zz��	��Z��r��@WMja�7���u13�Ys��=sF��-Zۜ]^�C�j�ē:��������C��s��X�Q�RM�ٲ�eKFE�aFDpp�����{j=��9�M~���s�C�p���i���&o�S��l}ϒ��У�V2�{Ƣ����E�)�$+����m����K_鄥GP��Ulx�:Uz7�o�V��Z���:Y�3s��{��Lޠ@��2�\�}�f �F�
��F�?.�����z�ď��-3������8�#�a9׸R����ðB¸	&��
�3�X~��/���
��/?��(�Z�D`���lo ��)�u��y��Q�H�-!5�jNaN��M�"c�GK0�_�f��z;X*k~,�V�=Ks�c�GژpT`�j�N���%h��8f�7�H뵫���1s�Åʑ�V�^50b�7ld0Ҹ��>���`͕Q��p�ӾϦ�ޓg�^�K�� ������vc~*��'�
dM��SC�ba�`-�Td�3e���%�Ial��0��v�a�����mFr9 +-~9Ā�*�3�fc9T4��n��x4(O���B>1[)v�OϷ��8옊�B\�"<�|���'t�Ž.K�n���/�.����ͱzu�����S��c��ə�;$�������<@�v��5�rf��?���+hp�����j2p/C�T_�NW���x0��L<ͩ.�8B������ZW��/��=�	q��A�>M='K����6&�'�����)HbuqMq�k�ϡN[*�:ၒ�[jU|.�k���x*�5$���h��E�Ƈ�έ�أ��rT�����Zk�Ѫ,�zۙ޾�k��Y,x�qN�0���>M�[|��;��W�j��
ez��a�XC}�-��:��R?p���y�o�M��U-���
������ij����y�Vf�D2�W��V^���*�hF>1��G����ə�C��l+8ij�7����x)����(�� 3b�Uˇ�~��5}Q���R8����`D�`�\�|Vu!���/h6�d�X,�Fʚ���Ă�<���*�6kp��6\%.�՟=cP���#++�V���#���u���M|Ԃ0� ��e6�T�`,u1��%*��g�"�6Z}DR�9���ί�2Tl ��m"����
���N����J��� L.4��\(�ȩ8Hш��eZ&��ŧ�a���/l�����4�lO��r��r��L&�i�}�`�X����6ndq�/Ԩ��t��?wǮ�%	�����r�M�QFoR �/Sd�[�����5)�27K~�� +%:r+���6�L�3��[T�7t�7h0��%�8�K�%.lC�X�$#�#ba�̈9lz-�0�ݹ1�?�p���e�Z8W<��r2�&� 1"�p��x	�=:�"�#ֈ`�~/������a��oÏ��z�G��:jʬ�!+��	=�|�%g״�+����4� ��hP�=s�J:4�ʇ{�g�������㷍�B���F���vK��+dk^Բ��+�	���r�N�F����Ær�"��MHh�1s�Θ�R�G�T��Ӄ޺�װ�W�0ۯ��C&�A�Q�iτ�8XʌS�7�+��A�M^�t��$j�jKQb_���g�\�)�<�}3�=;�,�����f�^GK���� fw�C B����J�Ox} ����!����~��o[}�o݊Dn��ߦ�LA�I���?)�ܽ�lYBPB�HE㑿��@l����m��^G��d�(��M�3��&���3���ېBS\�B�lɏڏO��Ȟo��;�� ����O�&J��*%��������I Ǚ	�l�uf	����ү�l�1Z:��;Ef�/��"�m��ڀ�j�V��5�Yr��"�{!�:�Mn���n��Rs�zV�}GJ,v酜��CK%9{!j�
��Ј�ME�AI�B��Ε��|+'O 8]L���yg�=B(�����a����0����,)q<�I?� �̓֞�$=��WwJu�;��(U Hdg�@w[Vv��A�^H	zm%�$�8���sC���)#����X#˔�k�|pB�7\*
+�X�-��
f�y����J�C�]L��j���������\�0k�3�M���zO	���D�n����e�N\3S5t��a�$UF@fu��a�:dJ��"�@W��j��ڔ%�HnA�l��4!�<�q�=sp��26� �ڗR���B�v��Y�O��� ���8VM;':�\�I�!=��ZN>3-=]PZ��5e'�Qq������j$�0����*�BP/��Y��y�{��-�s���M��,|a=	r��ߗ�о�
��\���;.����6<8H�%����� -�.84f�g��'#�=�G��`dL��[�С]��bW��F�ͩݎ�.�-"ʲ�c�����<�[/Rຶ3�@����*7-z��E�cVَ����ā�fj)Ů:`i�)�dҔ��3�q_��}nF�EF�rF���a����'7
�F8���$�[��C��X��N��p2!¤n?��urS��N�� Ѯ)kjG��X?�C���S�Y˧��v�#I��?,�]��ҦJ�fR�_N�pL�u b��I�`�bX�a$���q҅+�O�y�*8VI�T;��ϡ\����G;�_6���7��uCD���6ʄ-��\�7c]�l�3�����@&N.�~W���H@,�!�3^�y�L�Q��W�����D�F�wH����
j��uz,�چ��k/
X���}@��.������Hp�n����ak r������
s��ة�X-<6��c���I�s�X�FV횙Jޚ�n�F;�i�T�aw;i+�'���m�?�f:��CgI��č�֘�w#���W�C��,N�d-5�	\57�YI�	�O�g�3�؊kM�+�X�#�e��Ί���c�U�V����\��FgMN|����D����Z�<44xK��npE)ݡT�F��Y��#���[�Z��:��g\F���Uz _�Ӛ"J|�d�S�'|�ژL�N�3eaH�F����a˭p�[o����mY� ��ϊ	��v����q]=�pԒ�������*v�T�ѡ�����5Lk���\{����o�/��}��5���r�rڨN��_�C����^��8�u��Q���LMg���qd�c5<m]�rõB��� �V�`j�[m'�~	�46�G蕸�ୋg6<�N�5$�2p�lT8㧋�&�0����V*}T�j,Eq\�|��b(u�,+��%,�ЀJ�&���&�\��.o�!y$"W��ח&��K3�:�l��vj�x��������P�VO!LD�%���B���H�G�O]�T\��Z��{� ��x��;�����<c�
���>�k���F�/B[6�ȴ�%:\�6��aq���ܓC>�f�Z�o.tr���|n�#l�����A� O�����'�Bx `E�
�n$�vI����8��H=��!v�]��C}t��h�]��	fH�y�� +�M�"A��vC�"�kZ��D� ,�wy���x�Q�B���!m���������5bd_��m���D�Ċ�7tpR����,��̱6��~���jt��i� ���(��9գ60�3��h�7%:ws�iK��]�p����@,'��Tkd[7��?&���k�Y���y��#�T��BdE�9�{%4+��/ 3�
�,�%��b�NC�0�f�[��4*᪩�J|�<xjyȼ ��#�]U<��O�ڻ|�gD��z[��kJ��Rd8�]�o�V��{���`09��4��+��R�PW��K(�8x/8xM|�|:��C�&BFgƥ���w�����t��j8��g��Я����ՒFJ��i�T�~��N��?��W�-�g�.���f����{"�7 t�qm�r��J�^�mzb&o��F���
c�k�s��F��ҩ��㼗o"I`v)~� �	oiW���1���ީk���O�@
�,�%MH�C���8|�;f=
�KL����k��#�����X��x��@2A^��f�?�D��ڦW�د�A-E��3$�����&�X�~X`�b�z6ߊ�	�:�~xs�{͓!_�U�q��}N��g�M�K��
����עv4�,��~B���iz,�Hx�7�w��d�j$���F���PZ۵�y<�4#V���
(R5{�'�_A��.Ftw�������~Al�n�zS�T,��z�_T�C-�br�&��;w�U��OWc.M*��ŽM�ktW�}.�f�AW�ө��ed���s����B��Za/���|p�Ǯ^�e�g�9՞�	���_�َ�y�o7��aJ����B
QW�>+��TKW��2�Чf(��
B�|�w�_���$b7RK��(��~�3���厯@)k�b�q7�=aq�������4�򯣞������=&8ؖd?c��I��4>�́(6B�&�����9x��h��tz�K�<�
rۻXy,;J�j\�;��nSD�p�xr��x~�n���B��e�m@�.Ç���y_/D��͙�+un�^:��=Wu���,L�k�j�kg-�y�4&������*�Mw8�D)3��/����c�K��K)�E���i1�qϒn�����!�����:f�B{w,%��6��D=X�>���=�y���|	������@	���JNk-�9l�[l��SX.�� f��}�m2tn��;p�\��Se3��0�]����m\�-V}�Q0�yV��Զj�O��Cf^�,�<�7�G�J�s�����>D��AF,"�t)����T��) $�i���z���1�E,3�➿6�v�%Cd��q����V�7M�G#��U!Ժ�S�#D��_���<1	Cΰ�3[��Rނ�zV����*����D7;C�������`��!4w��������К�01��3F��ZA��H�� :����n�j��S������p�)�R��B�q�ܾ��.�<y�J�.�QPn�҅2�yt,�8����.Vs'  G(�v�]�����X����Ա��t{GgGݩb����d�Ǡ��P�qN�Ξf�D�}��ʗ>p�⤕S�͌P�����Μ�>�;���[7��I�{�����5��o��pϯ���SA�"���Q���ʲ��8�i�l�!)LI���O�[*��]Yy�-.��7=��WI3F�-%�D��%��	?KeF��h���p��T�u�U��<�������м��.K��=����w
݃uM=�ѥ#A�^��	��ۋ<9q\Q��(�e�+ ]�8�Yf��9,����R��6�Aw<�w�̧���\�l��nw�}o-��w�q�4 ���Δ�4����Ұls�R��}�X�g �}f��D���!��rd-c܋��� l��75���Wt���v�\^����t(������N|?Nj�Й	Y"����5�;eyhw�]`��ͱ� ���M�k)�3�y��U�
*Is�����#�*m��H�%��<�FkL$a��m���~A��{�\�a�RGK��k��YP'Hdw����]�c���(�����)�W�#�j���ֺž�����{�,hx�������ÕJ�\N�C�>�h��~���|/���?O+��D��g�A������(ķm�>�=�ޮ��+q�B��Gպ$B��Ҧ�{�ǟ��$��6���^E��V)��mA�w���6����%���ߜU� ��i�����i���WW�fpbn,|� iv��;���t��Qd�)��ͺM�a��ӄIȏ�&Y�\+����l�^(�Č����|,e�yn�5�`m��-�Pߴ�~k��y��"�
6�A����gi�TG`=�󢻊ȆP#y�=�3�S�?��P��t`9��h<���Z_��ZdrA?��)y��8O����]9<�����ܕ�ag��y?��y�RL��*H���=
��ť�8��!��)"�D\H��G�(%���_��
�B�K�N�����ɩ��dM<d����}*X��)���oM�����B�2� ��%~9I���D-�Yo�!l)�B�Rʵ��6�--�س�� >���,w=��ظ�$��Xh��������
�������i�4�q#�VSi��I%�5�ŞNG6*��Z�_G}&��Mūf#e�l`8��`��|�]i^B�!���"�ۯ�,��� ��������0���=*����q�cv'p#� ��|	[z��p��?lw	E�;�&���m.���b�h�5�x�t���=3y<?�=�f-������ى���;�UH�0U�
��0#����c�	�7���8rA�(�"����^\U�v�(�Wt�Dbrir��2@��l �q�� é&2x-��Z}��{D��ΔT7X- Иa\��>��	�M�f��Q�C���O:��N�J(s���[433��l�xb�(��3���2$��\2GA`���eZ�����R�H�
��8���i��٪>���������I�N����$H[�����yU�v��/P���C��Q�Y��Ҿ�\���e$�r���&6���0!a����'�{�XΦ� �^0
,H��R�
�8[��x�Wn;۲\��4$���@/>�֎��[*�3�).g���(�+Q�pg�2Vuw����dV(c�q33��!�y��"��Brl��k.��14t8_=�q4��<7����h�J������)׮j�و������P�'*�"/�s��!A�0�1�U�L<��Y*�0�B���}ݳ�Q^�I�y;�S�ρ���r|����k7���t>�$�v�c2JL�'�c�^"B�i{<���'<'!���t2�yv��|CS����P*��/5�'cӹ��%�9ɚ؈�{��F�::�/l)�H�-�{�8tk�H�sC�;F[t�R��,l�U:J���`���ۄ=D�)����W[І� ��׽
���� ����d� ���Ƌ��xYG_2dP�)γ�P �YX�Ǯn�:�����3OGq1τ%4B�-)���j���f��ᏢߋN��e�2"A�p��j�����wUBc�T�j�c��VgZB�wk��J�i.JY�X,��U�?�my��ҥOX�ה��d-O��\�|p�hd�N#����g1L�V� �W\G�p��K`��l����笳ăO�l�;���q�w�X"��M�����d��¶XH�����H6��[x���߮h�Ps
��ҼHr(���-U�����ĺ��Z���RV���b��~M2�o!,,���� o���r���hg�����˒쪁L���Ƣe�����7BO'�[�.���1%���U�@f<����9�˔�R�h�+���#�N.KsKe�O\h��y1�[����4����Y_C�����J��|K����.{jv@�!���c��-޽�̭]_��Áj�DiP=_���"��P%�0@���s:Ȏ]���0��)�:T�ɳ��P�g3����2ȳ�wi1�S,����`��U��e,�߼Lh~q���I�39)w���!�tQ-`I�-�𘹍�}�@���/��Wɶ�U\�G��6U�<�V,�Yj�#vGS��Cg�={H���'A$���t?��}�oj�ly[�v����ޔ?T��{Z�o�%�L�6�Yv���(U�M�	�; i����0��E��7t��m �n�=E�tE�]��h��E-�dlSqh[�	d:�w*���&��s�҇f& R��̿ٶ����c�$uT��,$9�/^Vf��ȉ�IOd*�퇡ps�|Bʽ� (\^�Thh�� ���6��x�P-�'���4�鄌*,U4=]v$fW���]��]�b��b��,��f"��g�"V��ZȤ��&C��xǸE���x�<V0��wl�ҕgw�=���=?:S�^'���[bv{�-�#T9��%��hУj�H_'d���##�q��"R��]���)[���훸���L�}	M��\0����GՓ4CRA�C4.���FZB1)'� q�����@I&Ƃ�j؊}��$�&R%��z�W��`-bC�x��m ��>ޝ ��0g��o�7�KI����q�s����3��1�tܷ��|���F�����
���^��byc�~���D?���.��i�� �ϥ]�O�5~:O}���4�Z�*�ޑ������
�b�Yf=�29�{�l�(��M2Z	ts�K�^Z�G���TreUء���C�Y̔�?Ӂ�7ܐd)1�&��1�\�2b�~.Kˆy�T��9����5�8?H�鬴$�e}��|"]M���D��6�f��	��巄c�sGQVǵ?��$�g�/D�!?���c�}�:L����T1uyp�9�"��P���^�s{q2�0��ɮ��6>����E��ԝ��ǿ�-�M��~o\ದ�ktN�vE�<�&�9D�p\kA�DKrϸL��s����?�>��ʲ6Wc���;Q!��z
h�i%��:�gECχ�����edE��G:�AZ�cM���"l\���Dv++2��:�&�����s_��E��
f�o� ��}�)S���V=M��P'��K����4-���n�X���(�N@���Q/►�����c�Lj)Z^!��x\:a�U9�''zq�&��DYT`ǎ�Ӂ�����r�[;ڏ�t�Ƭ��^����!���:񸺸Dp�$%��@�|�{�:��x�rO8L4�*&f��,������cp���E{�5"/t��7���H��l��m�'��Xn��7N�7k��ح%����ra~|(��:�5�f��_N[MI/?15g��ڒ�i���1����
HATԗ�*:�iø���i����?�vC�Ϭ2VI�HZ�OP��c%�F5\lm�DX`im��JD�F}�ٙT4�L}�Y��vv@U�jN��}�|F���+7�3·���+�o�1g��:�*�gey� ��@d$��n��s0e>
���\����M�����uv i�������*���Ƞp�I�%e��^��"��3Q���R_�� G�}(p�U�'��O��{=�ڏ�Q�+":����A�}8:f��70��NT[n��ր���J�M[(�p|�->!�i���A��ӊV�S"G���4�#�Z1��yg��O��B%�>Z�1�V,n�utA��G�
S�k [m�Z[��l_�������)�<$j/��0D���D�| L�\��
Hc�[	V;�u��D+�p|�����Y��TEW\���+��5z���/��Z��1h=���rϢ�_'}�_��Z��xD���e]��l���ț�}|��=̧����������I�)Zq����ͳ��T��gNDsj���Ǭ[ٿK�!Ty͑Chп���㟟9E\�x%�?Nn�9U��d��A��T�������Y,�8�S�w��P�rE��fX�k�oS@Yv��N��w��ӔC�
��B(�I�+~X=����i��>ֲÐ���;b��3���;H?��ҳ���rց�u��#�	��j������Q����)�r�:´2v�����ؿp!��?�"-�2���u,܈���ir�8��S@��I@�B2D�c�Z@�g^$�ե����O`0�Y,�P����v�l c��S�+�1y�N;u#*F�ֽ
|Y�Y%L~~	��X9"�V��w�CBd���Bn5��ix���~T�XsxO�V�kSZ��U�saҟR�g8��EJ`o &�p��lZ���N���pMR��~�Pi>w�!M3�_'SFB�e��W�Q7ӳ �Y(����+��n�_��Mƣ�K� ��h��x� Q��r�2�^���9��ou�5�RC4k:St�S�16"=��)V�J} ��A6�3������8�U�c�6�P�ǭ�ϸyb9H2s��UرqD�7������E��V�83��t���8�?؄H�U$���u|�cTy�������&��e���a�|�#*3w���o�( ^J��>}�0����r�Y����k�1Hleb�xg��Y!�B��� G]?�.��>��vY}��\-K�����1��*�iBo~rT���s�7�HD�KD���I;~��b��\��{�b�)j�n��V��I���Ǧ������]�Z<�������l�T]ł���=���ۮm���A�w��/5�'�N��!I��Pbo���}�p�Η7n�N��g����ũ����(밿��� l�0���24�߯��x�b��C� ��H�[@7�~��EFb+�e�5#�D��yk�)Q���jЇ�6�e�Qw���Vz���r�����C�
s��{��9�#�E��[��ڣ����Y�	d�,���U��ū�1�F��=�A�����'ZrR-�T,½]ȕ��ɜo�'�U�>8yk��Z�*��	��	�~��$�.0l�Q�v��6�o��W�>�Bc��b�8v_�i�T����ը��ܐbZS.��#���`M�"U��l,��)m���T�������gv��2��86	�N�QM����F�1*o������FI�vy�PҐx��n���8uj���!���ۂv������u�ٶ�_��e	ER�>:g������x Uܮ�����[�C*qr� 41������a� �\`R�ܝ(3�7��a%,[�<p�ߎ�Ϡ#�v6 ��kG)���F�!ҹ�f��뛜�+�[#��
��FFS�z��3Z6�y@�D�I$(��R��!.?{D��v���룠���.�yr��ϵ�Ѫ~��`AΦ6\ b�k��X���R�&?'�Q"\QvS{C*C�e��Vx���L�Q���%)��4�B�G,KY_E��l��^s"Ԑ�u�D�/�����^{ �7 ���K=!�^$�6�t� +��##(֕v"�R�]�?�J.����N]��:�}e�,ܿzrnaY�#;�6�R�����~E����<�E��U��2��A.����3�K�����RNFF(+RW-��o%�U��e��;�I`����M9�S��P��fE(����ہA��cF{X�@��%9S��� ���ig�D�΃�Z���Z��~
4m����O����H�V�}菓 :��$ŏ�-ݝ�ۑ+7[ɥ��1��(� �9Ը7c��)}�V��C���7�q����%}����9���'e�*}��#N;8�tw�W(���#[���`��i�pd�i�xt�%�bC�����NE�3��M��;ʃp��%4�[�mz%x��-{L�����d_�9!��ދdw߿��7R,"�\AC'$q��
��V<��d���q�� a��a��������@:@��v�/��j�La�т�7�����J/E�>�G�s��� *�1$e�Gg"���>|(��N�� ��W��0H��{��^��ș3�s{���\�/jJ�WN�Zd�?�w��M���sޜsR�=�EY��[�6ۆ��)	H��_�p����$�w�q`��T���6����b�{�pGcJ=%�^6Ⱥ~5�4�ǐM~DaC�:YQ"���nU1u�v�'�A�������t��^?�����QcdW+�C��v��Y������lP�������.(��h�K�ǅ@U���t�q�N���U8jv����x	��F�hRnd6��SÊ��N�
aS��)�n+�����V�R�+`Qy�oI،����F
��{���m|��ZE�
��T�/+�j�����/��2P�{%�;�UQ[0B�g���#j�ꋆ�rƱ���������5���/�^����6��τ��~f�DZ�twF�P7J��D������~��u俧��ږ��f����ԕ|wfa�w	�<���liq�d��ʵ*'�)$D��b������=|�=$/�狞���P��	*��YWH��vX�\Y���Vd�{�!�,=6����u��T� 
BC�B�ÊyP�����R�O�~"�4�<?UY�*Q�ΐ�7�T^�~x����W�q_؟0-���{��xU�-�,��6��L+�(����*�]DR��M�*�]�|-L�~�m��+���ڑa��&Ͼ�}�
�JM	z{�%ꂴPx��+�����BeC5�,@���H#�p�E�����C��������)3���h���d�
#r� ���"�~�@��W	��ھp��7���ѯ�^���.�:H(���HYI=z�����o�h�"�	�#��_%Ǘ��b�H�{G-r�J�6-FS�Ɓ��h7��`���^�����ho������'��~6�':%�<Q�E��Ƕ�<zO�j�C�x`�.�o�V�?�)�)ֲK��SР����J���d\���P���1��?�dK�4B6���x�؉�#�u��͌&㵽�r��O��� @g�P����%��IF���9:˲-��KH#���ޅ�,�yiݟ����������#�uj-���@Z�Ns�$D_���
�:|��` !������]lV�4
���B��L��	�ؘ��4��X��mp��qp��ª�V�\�`.7`.$�#v�@C��숹��{`�ٔ[ޥ��@��O�H���P��^
����R���)�|�?`7�Ï\L̷{o6VsO*��;,NV��[4���=o�< �!oe�)�'��.N��\�������)��kz���ߡZ~2�G��j;��Tt7�]|<4$���~ rlW��O=D)S���/ld�vwR�'���ͯ�b̴�J��3�IF 2�'F�"ߧ)Ts�����(:J�u.`�v��xu��2�4��
�r�2�p8ޣQ�(`�In��s&��m8({�v��ZR?TV|�Z�[��i��tk0�*j �����_G��'yY�\Bc���i���M����>Bp<��-�mT�Y����m%�a���q�N��L��<�7d!D{��N;��x�HJo`��m�~���G���t��|��"k��vcQ�N�6e?K�J���Ħ�1_�y����8������Ȟ��ɤ/E(�z�e�{����3�����G��[b�ʐy#��t'�D��
�� dNէ��ѹ��j�E�M´�ِP���n�ZT�����w�:A����j鍾<=�L�	�i�\S+�,Q¹���WBm�j��g����̞�2��{d;'��9�����W�m��I�8|8���na���sr ��"!IAm�s�5���;��μ'����^daM��ͦ�h�Z�[x�Њ`�`«*��� 4Nf �FU��8+�%�ܴ�xa�OS1�*U{nw�۔�{8�{#���B~Mb�ܿݸ	� �y5"C��k����w���j_��:_)�� ��|���r\���Y�,���D, �������:��������keBG���x�J��8@��5(B2M���b����kԉ:ݝa�-V�CAq�s���/Oqy-cw�*G ���������i>�`B�]�؆=�Q��p��j�DSRO��b- �*���>ƽhBF6���͟20n���5��4.���z�نpNTA����Fa�T����opK����˞��5��gѦؚ��9�WA���xQݦo,��6W� �4�F�oښ�0�&ŽǏ�k�`|�3':䠾���@׏�l-1�����P�瞕���m����g)>1��W�����!��I6���r DL?��ȸ�l�����&�A�Bu
��7�JI!W��_f�>\a�kX�B�sW�vT����$T�;E���cM8}6�����[�[O����}����i�S/����l,��]������c�K��"D.B����W��_�O���VT� -�ژ_�IN��;�)��5�ܗ�[�e\�SԎ?�����r�]��BI���X����0�A�7�`�/��XV+�×6���c�[P���(a��c ��C0�O�|j�P���.Z���*��r�����y�\"^�*��*P��jE]��Q��}WL��țZ����kJ���l<Pө�_x��A��y�Pڡ����p����Y�CZ�T����/+������|��\)/�Z���D��-��^cX �a�������kQ7�-ߏ�c(���k�I�Ho8�.c���9=ǿx���v$�޷���BΨ�Ѽ��h��nz�Mn347�|o^�Yw�^�g�~���zZ�tRj�oJzJ��\7�*S*�a��c��<�|�b�w��^G�ж�	$|����~Ʊ]i@�9��M{	(��d�7����K��*������m
FN�o�����w����jz��Y��zQ{��a�Q��f�UE�,�Ȃ���̉�FO�$8_�θP���*Ldu%~��+���)�.Ȏ>�
<=���Mk��Q���Nl�yhqǑ���)V4	K�H��9��J�/��!Cb����P�r��tos�Ho:��v�O��iN����:�a|�i�}u��cN�s�g~Z�?â2�:*�W�4����3�A�c^�Ͼ�i�ud���=e��y��I  T-y�\+�R���qjdg��^��m�8l�c4~��=4gd���m"5|\�8ISM��(���T�r��9����B�����(��5�zr1�.�x V��Ƨh}0��q|��30������NK�!`Z�Y���}�M��-��M�G�q�^X4�T��O�h��<t�����[�V�Q��e�Y_<>�йA_��vϜ�v���D���$ >Խ�s�'U@�[ZA�J�w`���}���U�2s>��)���tg?p��?/C:���@��q"�����l�
W�����h�"��zo����#h��/�H�{"��axl+�Yg�4A ��i�;���g�G���a>L�,_��� ��L�ÛU=i�Hs`�q��p���PDV1�E�&��z}_B�ht.����yy�c������v_��G��N��:|q8�MiRxd��}"��5{psF���,<Bz]��ܝ%�2��W��|�.[������Fw��g�r�CBq����邦	��}���ANϸ�q���� �����j|�$p����#I3�A�.�Jt���zvTQ��Թ��Ŷ�?�K����L&"�rh#�t���b� �|�YG�7Z��!eu��`H+Ǭ.�0�]?-���kN��3ۥ%���ϼ�L|yD�j>$�=�f���{�#��+O�%׍FƢ����c!(��ͷ���X��=/��Y�I\.���r��;W^�v~��p���)Pa������2�r�S ���(�\��7I�d^����t��$�x�u?A�N�JH"�q��S9ˎ����'���Oh�=x��!q���VyiP���/�9l9o�m��B9
oA<�6����M̞�������I�&K֤�����H�mK�T����YW���\9͠�։���R���N-��:z(�~�d�����2��a@n��i%.��f��Me$���6�%��V�Y��Ao	�4��K�w7ؗ��1��T�}��|�zh╢��y�?�̯��U&��8r�4+F�.�����:)����U�m��Z��'!CD=��疡N�o�L�|���c�����Y#>A��T��5^�ORV��I�
���e������r���9�����V� �wr.����+G��f)>����D�8C�6���$������T����� ��\+Ci}�k�qjs-�x�w6��w�Z8��@�GF[�,j@�N`�>Z��<}�.��MZ�R�'Fΰf��WJR��~�IpE����uF��	�=vJ�j�J�#��������kj[K�Н� ��'ݮT��-����s��N��ٻ��
de��p�T��KW����1�PU=���M*���E �Ͱ��sd�B�_f�m�rY�n|�n�?�C(E� P��i.	3b�5ћ��&H�M_�v��uy�_opJP!��7T j�aqF���(�^G�J��i�|m��ؿ���
/T��~f7Z�e]�M���R��o��?�k�jʠ'�[7�E���1t�o4l� ��t��*�f~9g<$�`-��{�>� �8j�N�L���^�yZLN��߫k��%�#B���Ɲ/[k���Ʀ[iB'��Z9c]�Ft�/�s}*�	rK�T��E̾95T%�����+�M���C�i/�
~f{�.p��,� �P2��о���g@��J�e:cEĦ���G��2#l�g��:� )���!�xe>�v���m�$}����n�B��\;B��99:ʍ$UI��TF����T�Aߣ��ֈ�i��,��־+�Ģn�ȁad;�ǣ/d�~A�

>v��=��攮7��䊚�I�"��֋�r�qTG�i���J������]�A�:�#
(�]9�:��u�(�S��s{~�Rf^<�F̂a�\g�6�Q�)��+I�����r��^�a��.V=@��?�GU��.�/V��`�*@d�⮩���C��׎4��K[��DC�bԢdヒԎ�5���6���n���S��v+��n7��)�� �i�
�P��T��k����fKm7i� X��tr�p!�z�=��
~�0��"�,�Ӗ�u5v����\��އ Cq)!0�qi�8����آ@2ӫ��'"��gq<]{�|��*e��/���e;r4f���8[�\�L5QW)����j���� �l�����CT����/����1"u�m��.Bˎ���?�>c�W��j��~n^aV���-5�/Q��PdfL��Pa��\�A�ޕ��~6V]�>�\#�V? �� �_�J�A9E�c���=��-���	ⰼM��1vz;q
�
���y�g����X�U�NAK�L��!��%��ȓ�[6<������r+�A:�V�w��P�0�51ݦ�{BK]��Tf��N��!�
�Ť\���)�o
'�3�b��;R�ndG�:�e�����~IU�8U���D�XgҚ�<�"���^�#:Ƽj���a�kʦ�)��B�w%����}���t&5s�0cG��Y �	�O�C�fi�57�ݎyiJ�n�򚽧���8��� 
%�k?��y��n0G��e�p7Q2e�膨EG��T��(�:���) UQ(Z�O��P��,��Dnυ=�a�:i�����$j��F�ݓǨ�C��:;�>E!q���x�o�By�7toiρ��[?#+�&����iq�a�Ib��H�!�гFi1C��15a=���#�-3y+�$����p�*F��z��ٝ�a|L�����0�h[_��b��j&���i%V�x��xlvѩ���������������[}����V�|H���.������~�B� ���/B�;*��n�H�tAK"I���ԟ�� Ǽ�,8*Q�n꯴�U&t��t�箶UxB��S+yW���tL�PMr���[�G�`=3^�FR�������i��9@^
r�p��̞��3���>�N�
�C���{.9e"�\�LhBP�Z��"�P
D2�M[J��|��d�����Y��Z[B�!P%�]$��$\��ᙻ�h��Ŕ�[7=��lw钬���!8Pp*m�%,
`��Wĩ�#f���}�T���ѧ�mi��.�u�G��C����J]��j5���Ja�Y��6R(7��e�"�'A_]���ì��(���'����q!H��'���0�L���>���A|�|����R��0��n� гt;��I7<+���P�r=��xW3g�r���G�?	V��'-�A�s6]�4�����l�.&#�N��sZ�+N)d4;���^�HYӳq�i�*"���_�R^΋&���I���QC���{\%�(����kN��t.�c)e�K�j4�:=F/D�=��4R�J��V�ȘD͑�9�x����K�'��G��gE�򫔸�	E�`<��;������76wt�g��/�D1<3p���7�S�2{V+jh�d�L�?�)�a/Sm���w�u��SWMe/����C���L���Я��Tܪzl��[�2���at���ǐ�*Mfqq%UM�P��f3}�V�>x4��#c���S��G�>���}(a=J�w���_is�(M��<Ѹ�&c�V\�?^r�}0&Y���.WK���A�Z�J!����)��
n�>��H�����|XH��J��Q�M�����-uqK,�^Щ,�JK����KTExx�A�y?�_H%	�3����Mo���b�RǬbbǳ�0ъƍ\�ʆ[��ac��{�=���yYRn��,0K3>K��)%8u`������r%exT5������_�E���mX�R5�g�T��NU�8�@ݩ��#Ճ��2�yP5��G ��r�o	�dTd�բ:�Y����%3h�OzލP�2Ʋ�B��Z9	�@�0{�nsR���k�|9aBj�2M>am���:v�;.<"�8J�7�k��}��?�M���W�4e�x���4j��A���Ί��ސ3q%�P�G�3\�s�p
<�M�[F��>mO*�U�}R�����S�"0����ȸh.��,���g��\�⎂1t��d� �=ݣ��dֺ�]�������=�Ϫ�h4�(�>uuS���0�~w9���5���b:is���ɝh�L�A%;J�ӗ��7��͜�y�)�=���#�����M�I�s�<'BE���(ɮd�6��3�����e�Y3\������������9$N )ɭ�*�[if�*D�	|W�a�����,dj�������� �$�9��x5&UN���S�D���qa�|�������_�T�����"#)h�V��D���l����$�BH�Z�,�F���U�2�z��v�S4�y���}- 彇#mO3�Y�zV���A�s\���[ܪH��\g�ܑA^K�¾����V�!�RhI��U2Ŵ���H#�i|k��z3�G_m�rۤ�v�uSؕ�8�YN[�u�,������ip#���8�бB��N_I�Qy�&�h�R�����m���'n�mÚ���֓C�T(/O��	�rq�@g:�x+�˨\ܵTe�Lk��(}�Hz��
T?}MQ}_Xd�u�!�A4%N��JM�7Z��Z�,dC���<xQ����:�^�0�U��JEd퇅�S��0GG��y��K��@;�\�9Q~��N:����	~\�%��C$fn�blQ@oPE��]B> 
�ܗM+"Pn��)���QntG�q�w�-	�@��L�_H���N+�H�I'i)qJ�Y���S�EJZnL�rǒ}��((�㵗�K0����g�$��A�B�5��71bX�V��y2����[y:�h��ni�5d�}�����	���N���ʿ5gcճ�����9�W }�̭��n�-;�39�p�\a�|-��tXc��U������c�&_#f~!�,��ҙ����?Y^b�w�іſ��xT>D�G{����㓃Q�W�8O	���� �z�K�t����f��ݖbe�rE������
���+����6r�����F�_ ��
�s��a�P��#X-)��%�l����T�}p�WV���vb���m"�6@e�UWї�ԡx�!�{]�K�_ղ	S?�q�ɪ��9��Äx��҂6;$}QӤ�X���q�b�����L��8+T<�Ϫ-Pg6GuAj�u�}��T+V���?|4���2l�zu��0�k�
���]"bqC�ǩr(W��������Cf\HC�|5�P'�K�?K�\�L�W:$!|�]z}��6%�e��XU\m�.�֯FqR��}�h�!Vh�:��ٖZ,| Ios�Ѱl@I
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"��ڑOrdZ�h�? �sN��0���n�r�(����Nn�]fw��L��ہ ��m�~��E���Q���@]޵�Y<^Ȣ��6^��k�Rml���6d�S��?#�_���AxW�7J�*�6�tʺt�1萐��3���*�loq�KA^�ޑ�[�X���s�s�ɼ�1�O2����M���/~���m�5�w.�Ɣ��i3	&M��c�2�ղ��FgtZ�1^��>�;��qGߤ�2�>�mf\����s���w��|��xW���#J�g�Mc����������x��69��Exw^��O���e��rŰ��%A^�YO�}��u�{��:璼:ܺ v�7�w���x����	-�~� 5۵��"+)o��Ƃ�R�_!84���ͦrxWx�X�Bջ�A$A��П�T�)ˑ�G�_��Cɀi)"���"�guE��j� O��j��s���(}8�̲����
+�L�ʰ~����Go>{��zN��`0p��60>2�k�fF�)��A�� n��l7������}	=��4����[��q?�� #!���ND�5��z�f�&e�^10�io���	�T�@f(���=�<"|j$���]\�y��f�%Va�1U|�>�Yi�e��i�xpr�:}u�H�p�����,2�����ڄ�����p3=(�Q��	���Q�C����N��Ur�.. ]��j�M��� �g�5��X��d0��[��|h�"K�6����f|�����(`�% �M^Bv������Бʶ��!;����"��_�/��]�u���.��k{츸 9�˃Fğ%Vǩ�!��j[IS ���bf�� A`�ne ���/1�����O�!O�ص���f�3R��Q�akfĢw��A �V�Q���I���Ѐ2�(�<�t����H��\}2 d��j�(�[uIZg�ELjW(�pOaf�W�D��f8Ks�Oh+������d�%��[
�T��o�qM°A�T��佘���������;!ɋ����1�v7cg
��V��u�c���NI�&ъK9M������Fh@94E�p?)�Q冹5�o�F�ɚE���L��}�������N���ϥB/B�X�Y���播s�P������@V?������1~3;_V*��:׀���À��e�?�lץ�Lyk]���� \V/�x�h�~�'��>�Hi}�	v��"�W�NI��rU�x��I��i��I����1G~F��~���P�����C��-�,�>�=�.�N��9�(BLF�BLJ�CW?v���e��#��9	KZ�TK�<�y��jݶ�.�q��at!���Y��.u�8�*}`�d�Vn�ʸ?1�emM�/�e`�GɎ��%�HH���Y'7�--BB��kݤl)x���`ܾ�_�	og��iǃH;�V�aV}n3AhH�]��-Ip�-��K��eH@I[s���|Q������&"�Ȼ�.5���Y�x#�o�(�(�e��9�I_����u�L����>�g���L���e$�#��������r���C�y�d������3��w\t��V�Q#f��O7�n�/���N�ҷx�SP���F�Ăw�hWI�iۖ�k:M�e>\��!b
�r�`o�sk�ko�~�j��\7�� �7(�	�v�덗�6��&R�*r�4c>	�ѳ�K�
�	�
��$��'IA���|�����e2�>���5_N���	�W�_�N@�y�0���\D�ŸBp$�����f"o�vB۬ԢxEkV�qbHQd��[�oDQ�9�F�@r4�Q�K�E��G��}��F������\"wD�@-��s�����i�u%��t�k�5U˾`L-�y����|�h� 򬏝I>��"Tx̎_��L[�j��>�+���U:��lO~~^sc���|Эg�5x�Ef?`5��T��΁�59
m�d9�^i�-��!���R�AsF��U��r�l�?S:�f���C�ߗ�>���ShA�F:�O�B�H�O���}8up��JF>|�!�X��o���`�l�?�/�
���h|��4�ƃhV�J���I��2IG
/�u�S�<J�GbQ�犖o�ĳn)�b�:�pr�j��?�G���s��.�jih ��ݍM��V��>0�=E0Ri�{Z3�-�יD����知n"�3)q�k�猂ȹ����?������r�������l����
1"�s�D����ceQ���(8�S��}M{5�q�q�i`־ϯl�ra��{�S�v)!�ؖY�ϣ����L��.��ې�a,4�$��K��$���h5��z���V�v��m!@�i�D�vo���|�Z<�����CYR�dz�<k��"�D��?,�V#��X5�(deu;�ɰB�x=��<b��4����tk� ������v���(�Ҥ�`DM���d�A��DP���Otu�k���^}��yY�E��Q�iF�gkF��v���D�NQz��g�M���SR�ڀ�:c��G���v4+t�/�$�'�+�`vD2�i�����%"G���~8���YW����	����}��'�7gg��v5i��y��س̥ �����d�W/���D�Z�/V�42�'Y�,�o�l��d���ݖj_N���*	:��3��~)���°������\Ф^ޅ�/gj�j�=I��&)���/"�#�}]l��9���N1�Xy�ր�F�͊��XC�+�F��Ih";�`�J.ϱ�#��B���W���-!��q����MP�4��p��3P�2m�:��૯e�XH�'/�O9��b�޵��o��ö�{�3{ʇH�=�;piq�L,M��YMH�|ȣ&�E�O�(��^�8}�e|�ۑ�H�2�E�\l�t�,k����
�0��iGe%˞hh���/��,�G���oXgUlu`	_�|���0��Dw�"8Lxt/Vc(�z�10��G|�Oܱ�>�����i�n�(>���,�i�� �iU(��/5op��9�\a��ϫ �&Ϩ�8A?�oJ�3AgǴ�W.��B���8 ����ӊ��a}����I�W2�a�������k*�m�����$��Kӻ�u�)���}4d����s�<��S	�)�-���k�?�#�k��WК>I%�I���3� ��Le�e'�NF�Y�:yB2��r11��=Q(G�a����G�b���`�zǺB�r�d��>�ӣ#˔A�^'w���e{B�w���c��WT���dj���ҿ/���\�3�h��lf��2����I��&f�Ճ,u�%Ì�B�%�;� 9��`AІ��W=N�R5�_dh�K=�r�R�w�YZ&�F�c�=lD\�8N�ou~�f�뾪�"�~~��&q�U_��o߅�TD9�Q�z|���O�R��	�7��f��uA�$i(��t��(���!c��Zzf*s�-�f��jd'�m)uL�Z��b�Y/>7\^o�OE�B��N��fφz�^J�y@ ��;�IT��(<�<����.3��7v-(-�U1|5O��!q2E�E�6\#�ց�ex7T���m:�H�w�<$�&ǡqu��m.f�0;𾟅�%6����AR��9�z�9����O��/�0��g��V�;%�q; bn�B��ʩ����_=c�� ��D����=�<�&�u ��@��lA���A�e����"������Wbw ��)���&����q�
�K�������-���I~dǈ�$�5��K-Y�6Qz��t���L.5"鳝v`�w��@YC-��c�pc!S���Z,�ܠ��������09��n��/T��������)��fT�AϿ�)!8��J�>?a�����^E��HK�q���{N8ߨً�ӯ�
��!y�i�[e1	�p��8���9s�W.J�oK���F~�٬>��z�v��j[$H���gU8��N��%�0�tǸ�<��j���i|<7l�ؠE��!MS<G�j�گTA7�RශDe�e�������F��u(��ܾA���ʅL`V*��Qn���9�-	}|k%����N�R��<@�� h����=���E�S��xky���k2_��{�뉙�ќr 	5�ubl@��??�</JiS��rX�M��!�kׄ � ��)�C���8C��CE�*G���l���>�
K���V2�Y��W� ����G�~H��P �Ք�����x��W8�$e)O�����Gqj��?b��8m� ϯ���>�s޳�ӬI�,{�]`�ˈ�X_ �ð��=�+�P�.E]B��B������h4�*)o����~��J�ák�\�Q���8*�g�5�o��#��^���o�|��3��s=+-�>�+�%��ˌ��t�痨�@�����`�D,��s���S��g2��̃��Rv�M��A5�l�>�`2�� ����D�$'=B'(�!��xdD�wkԀ�8�Cj��w�#v��2έs��Wl����'y�q��앇I~T0K!@C�Y�޳���������Y���&�P���S�[�_|���2���|wB;��
H^��uzx�A(�m|�u�j�:�&=iJ^Mʬ�u'G^K��>����}��U���K>B�� 32V`)�_����2f���IG����"�H��3lZ�Zƒ�����t�"�\��	���A��_ـ�t67�C�\!b}Y=(z�<[����e�2�}�s��X����"���k/�����^�qK#9W�R0|>�})؋SH�w��*w���mOFz�7���oZ�
 �O"���%k��{d�?Gg�$D��$��TCo�u݁S������Vw��%�.;^z���O��`.�.K_x���]1�^F���	���3�X�فơ��ц�����w�	�r�ǛS�������邵�t��GL!��(/0�0�*�/������"��/c���[{������4-X]����﹞G�Ŵ$=��H�ƃS�/[$��ts��V�P����L�'�XJo��1����i��Zs�
�!@� �Y�P�I���I���U������� ��N5@�8�'n�6��izb�g��] 	��}���=J b�cU;S��x�u!Q+�=J�T��L�V~��dw������O�hr&�;�O�J|~���b�^��B;�wO�E�����ee�r�,�h�����0[k�^CN�(A�=�xH ��C|�J�f��Y��[Mr�Q<��Y�ةn��-�)��w�>NX��l�E�d�X^������,�:�,��g]�3�S�ُp�؁�ky���'[`�Y��� �[��������3��Wn"�C�4��1,��q��M#:v�fȀL-BX�ZΩ�'��yk,X�s��R�V��~#ݱMR�V>)V0�,���R�r1�|���F��J���5��U�u�2������}�y�V���^�'�}�����儲ņ�a�aPh�X���4Ǜ���!��[3d�*J��E�GS{(}V�
x>4D��"��.U��^��V�Y�y|�xr@�F����s�Y�bZF�Ά�d��kB���"T���<��Eo÷�E�p�����{�U�2�x��Hk�@��#��3�|�����heli������H�HF��[p��������e����&	�P��Hs^�H��'��}>e�9r_��M����X��b�%�S��M�����̅��"� y�B�P�M�=x ;�wr{t֑Q>��lmi�¡�~!�섿��$~fS��B������9�q��,�����>N P�r��'��^�t�@���j|ے�uڥ��9�g�Q q�����}Iv�Qn�[�ʱd����8Dl%	6\���(m��5�Iu�'����J����c�����ꢁ~��VG㿧�m��t}���F� Az\u]���솳�u_v���e���׎ܣw�`b��Q�7��"qgX��/~��̂�F���l�"�x�O�4v5�����Y��N����w�f5��%^3v��f�K����S&�7� �Ĝ*�j��q�����@�"n������H�J�������H��EY]7�ݐ���x�hv�Z�wߤ� }��tȔ|c��jtW��� X�yoQ	 ~[�A(�Ke����9Ē�NC�{?*��{
PU�M�X	�Y���ʸ�F�c��Q���.<]�6��z;�c�9Y�����ݸ<��e�mC������g�};G�V#NT�@����ً� ���S�v����\�T�A�uK�����6��l��,u�v���!�G�B��(=X�q/9ň�n�%皒��#斳U�9����J�6�Y������}���ED�Өx�p��s���/W:�2ۇϝ�!l-e��_��$�rt�M�o;Sj=T������
+�Q�=�p{�_c�9��>w� �¯o��I˲)܅�o�2��'�N��2
�c!�U��ϧ�0O���]*B��r0}`�;y���r'��)Fy��˯h5GD(���/3]9��-��V4������,~���t�s.C�M�J�'��Y����V.�krc�~4�� p�ߘ��� �����<#ug� �����F��W��F-z�>2�ӑ�yT^��̨��R���N)�*�[������5�w�$�8�?�D@f����B]�.�Ta�n���v/��kj���Ꟛ�w�1�d�0��!�s�{:ȠX�ܤ�����7��L��9K�Î&�=@9;��3��:�o�,���w����+�Xܶ��%�E��or���2��ƒUOu����n^���������l��G��*��۬��=���_&]����I1�y����l�q�V�R���r��4-2VU�x��I��<���]wMZ�ZMsf�iU'�Lx~&OU�Ћep��O�W�Cp���&�&�\.a�2v���2��.���H�^7W���g�y��Q����u��c^��Ma?�Mngtx�����P*_�囿�̟�X�쵝��Ծ�
e�)E�U�"۝�X��ã��@K���0.��S��i��
��1x��ګ��]~���~��nG��`m~��E�D�7����2�[��	���+�r�yWn���kh?{��ԓ��}�㩹�\>W�^����p5���Wk��fu�%(����[���;_��w�)�D��wS��D؆W}��K)�w�A��a�ꅔG׶�rY����&��7�TbI������ ��!٨1���������U�-��7�/n ؍e/�3Ѱ��p�Ep��(s
o�*���k(N�1�d\�~��p^h
�4?]�����DymVt���`����J5I��hP��D7̰�#.�ixGo�>��1R�)ťr���kf�n�Q*r��MB��LA 5D<-[ i�*(³�ͬlZ|Y�l�}��=��D���r�MT�J^�~O�8�Ol%m�>$�d���>������	T}�� ^����犆��P{B��5-���̮��3j`a������P��y��"n����ؗ���_(� �=�XT�rs��K��{�q�|��`�
X��p)xfV�e,pp/S�c�!,��q6Ն|[���� tB����M�l�d{�����~
Y��B��\2~�Y��R�����^�5������	)��ž�R��̹�]e�b��E�;�l6�[�V����Jp5��jqUP�� �a��/�����X�;;�vWj���=ץ�%�ѹk;I�׶�!,e3iѵ�unZ���nˮ����d�L�ޢ�L��`&�.�Rf���lluOuᤶ�v��*�"��������G��b��[�Ck���ޢg>P�Nq(�'��/�+�|����x4��� ��-�.��?��q&Z/��B���wY���ρ�08Ts�����PLƽ��ʇ�C��,'@+w��qhn��L����nf�oP\��f�?9���4m�]�X��Ek�v���L�!d��t&�!R�!1�O���p)JXz.�pU�W6�Ҙ�{���}Ġ�WF�B�J�J��<�Յk�$T,�����C*�����o�4x�.T�Ϧ�FX��Z�PAf`LA���gI���[�x#FӇ<6���H�h$�N�]@����O?	To^}��)L���7�r�ȅ4�L�k@3�k�O�q,�f���X�Ic��K��&� K�:A��׸Iw�5��#����,L?�Zd#�����;�{���<{�w����?B^��TDw��b���i���RY%�~(L`1uT�B�GUe�-��^���/�t+����:�E)��%�M�i�^��_e@��1��""l�"ϱ�Dѐ����k���b��
.�G #�G����e�I&
�ޮ�.T������:�����F�z2��<�S}/q�^3�+:��x	v�˙�y�j<���8��P<I�LڝO����<!��B�D-ر���;m�Z��M�Q��_���V�k���1��L	��C��J\�C�Aj	�m��#�*Z-%#�d�D�a�M&������FW�p'Jc���눕ˮ��$���Q C���H�Գ��p�4����=?�����$�MoN^�wݞ�?��E��||��n��g�dW���\����d��b�$�����O.��L F����*��'pJ�!Y\���Y���h��.��t�&�\� ot{;��m�8�5�#.�֑,6��sr0��8$T�r(������<ĻK��I�t�_{�2j�o�ڌ�����RHpʟc��d2xL�t
�7�����������p���Iv��z�zɒ���Σh�$��c��N=<�����]+��y#��G���z��te����a���yx���q�*�c6Te���;{�l'N�M��c�J��/�K�D4�Mj�?���c8��sS����uו��܏�L��L�ј^Sg�Q��b�/b?��u*���g���tD)٤b���.�o�f���d2�.��|�>��,���>��8�XN����:A��������t\>,x�4�{��)�����!oZ���T7��y`�}N����9��Br��NHD_z�h�FN�&��$��v�=�q�L܄���4�k�'�w�6�(E�V�� N�r*�����V�C�K�A��4}��^�8�0j+,�W����u�:�V,�v���ԉj�����I����)�j��㤸ƾ����GzKf���aėW7]�	��F+�8���f#�H7Y��pD�8H�=�4�$���]��LC�����P�-�=��W4�|%���F�6�ܧ�7���B'@��^T�v,GTbW�⬼��$�G�$���	-�H��I��&s�R��>ͷ�~�ѼSe�z�%����H��V��|�� cTiVne4�j6ù�R�����|~ґ)��E<�q���;�:�A�4�����#�A�m%XJj���v�����[4�̙�`�{���{������'�
N2A�
�Tv�sjImAc:��=��ckY�s�Jן~�i���2폖�(�>�V��0/����X�j�g��D?wa5�h�vj��&����k@�w��� ����z��y��4������P>��B� C�
+5
��'�=��y ���K-�W@q�T�Vw�gD����sހ�lo!y��׈��#�zʑ��0�F���b�'���ii���U=�%����wk&������/�=~�W�"�#Ձo�� ��[��bvGIK�C%��Y������xaQ@��ҟ6��X��0��!N��ы ��0D���57�7n,��D�= �o�Q��`����~�ϥ�e �7�{�0(S�4i��d�7  ��v����@+�0��WLإe��q����:%d���`7j�2p-�����mf�p�N��k{N"=��>�տ\w��b�W��������@%=��Sh�W�W�%4 � !�U��0N'�GS�LX�U\-?�3�C�5 Өb~&ț�&�kjv�;�o�>�(QJZ{�|KW+NR;`P��U�4q.t%��M��"b�4Q�V��]����n�|��xgy��n�����J��ZGI�S{���`�SWN'�?��*����6���Ыǘ�9�)��T�Y�)�Q#ՀM�c�Y�@B���bn��E��*e��ޞxV-3Iőv�u&���ߏ��y`��_��49��~,���J�0`���&��=��w�2�Cٞ'tI%̒�Y��W����W�]Ҟ�Y'h�Cw�j�U�bS��Ѓ]RY.LN�m_� �F�����J��DWz��w���*L�z��]_�S+Cε��<��|�.�**���	��R�6-m�$7΃� _uKk�dY�Ƒ�O��dq$���I��ΟE����V})�L�������W�~ޮB�λU��M�.��x"K�J�>�Z��Sd>7*=�޲�yn��rem��S�4C ����>t�a�,��h�N\��/�Młܨ�ق	���
|�qpxT����	S���(�)��G;�������Yk���r�ͻ�^����Z���P�z-pT�b8w$Q(Ԥ�Z�����w~�p�-���#�ϴp�wNSi&���o�#����㗝`ʓQ�E	V;���L�3����42T��'�y���|�,��#Νm|d�" ���N�$���q#\GJڢ�qvcƚpB�7�9��U�5���^ȵ�����@�Pt�Tϧ׹�RG�XD�}�}�{]5A=�<Ak��	��r_` &�][�ܢV��T�*��,!^H-o �bV��&b�C�bN5`�?�N�� �og�}h��.dq��B=�݀���Kt����BbR�T /��]�Ư�n�C'���	 ���ϑ%)��*.�:��Z( GB�@+��T�9(���9p`����-�NΦ��V��;��ݗ���I:P��+�߶�Ӱryʺ4V�%	�4��@J܀D�{"@H��T�:W ��@e�6:��$���!�E�B�N��$�|ٺ~K�\!��ڀЦȦv�}d�g�E�P#ʛ��4O"'��u�T��{�2G3��ǭ���{&���ʪ���̥���Zd�]x2w����Z�f��R��(KqY���V7U��YL7(ba��9�P��o��r�%� ��G]���>��ڐ}�	E����-�� �4H3�0�Z�oMa@�zխl��ɖ4<��3L�������mk[r�ҝ�If(cy�Y̍��ƽ�4bV�wy Sq�r�T?!���F�?�fX\��,g��C��,�2�]|�ﻊ�>��gOp�J�d����_�J	_yN���x2=%5�r�"�w��>�l��1���*g�A�Q9�u=�i���n�*��$�wy ��2-
�����VW��;��i�+	y�,B�o0�jQ�Զ��Y�m�t��M��HN�QM����K�Ŵ�r���y,�)2�{��������6;|����������aʷ�b��?���.�!=�����# x ״���a�?�8�|�,���6z�A�B;�|t)��"�'��D!�¨q|��j���0��N���g�`P������4D�_�PV�,�$=K+�������!t� ��⾨h�O����R��a�eЫ��j��B@o�Nh3H�7��6\W���km��/�E��)&J���zQ�b�:\ۺDS��.@L���L��|��~@�p��*�\���P��{}�tj�y��ƨ�r�ОoEEP�����x�]F�>��LU^d� �hX�'c���'M!�,��/�7���ץ��Jw8�'u:����{lQA��K;�(�n�<꤯�4D��t��Qj�f��u3�[.�/��y�
�]&D��AmΧ�6!c6��(9�;���)~�ʭ4��u�|kux��� d��5��:	\��B�-- �����;��7�;�@KYvr�)Cl�0N^&�o��T��Rns����X�ꑚ�э����o@��-?˚l�$[�	K�.4>���t�3y�"�d��7��/�����)�����	�%�jP�����C��%�@���W;)��t]s�݋�C6$��:�,��e���>t8.�����B��K� �� �p����$�-L����t2���s~M	���_��3ذ>�
����:\�ﭡ�f%���*��~�ШyU��r�}�M��[9wE,)��X収Y����6�[e��x�����t�v9{R�v�4Ih�����{w�Qoh~�}}17���?�_�Lυ־��<k�%�����j'���PL�K�h.�gf�������=��q��r6f2h"6&/_��+h�~L�}�nyVRL#�Xd�}rO�M-{�4��e*� C�H�Q\k���(>�-cr����?V�BjtF9���ab��b�O̋O�y�=x������<�@P�"�c�����x��<�)c�\���j)$!�8��dBJ9SR���H�q��@ͯ M�~�a�e�	��Q�`Y�n���,L��> ���~V� ԁ$?���@��2}��eʋ��s��������g4��v&�otL�^n
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���r c�Y�mI�1M�Adb�t,�i���ʂps"����1�BEp�e��mN�Iq)iv�������K�U��W�; hY����:Y�*�1�"#�.Я�&f)�MM�^�kt��F�&�/��u�Y܎�2�Q���#SL��s�Wl�Ȉ2�s�!����}��u�R�\#a�-����!�
mD!^}Zu���D��?�
Uí���6�sp��:���$
~��H�������e$�!^�0[�	-Ӊ�q6�Hm����^v{(�!�ֶ�|Q�^A����*Z��Jֽ��gI�t#����`�kT%(te֐��(��`�o��ҍܺ��׉O��	���]5:w�m�+Aj��E�������
+�sF����w�7ݘޮ��?/Õ��SՇbO��wf�Awt��_������"�O�c�l��|�n�J���@a��sY��� �q�4��mY?Ҿ&�4�w�o���@q4s֡�t,^7>��P�����!\��nl��'?�=Z`�łUS�v]��r�RTC@Д.�73�#Զf"�����|Dcx�ʆciLoݽ�(l���.^�͜�a�6��!-߼�cs����f<:�Z�4/���X,&�+�Jb�A}�cg�K5k�NL/.b�Q�"/����^@5�l��5��T���� ��N������t1,���哋������y�>R-)V/X�	Ð�������`�Τ㩾U:ȵ�֯����m�?b
\.�0Kd����_�N4��R-zp�=.�U��s��y��j��r�v�������@�9�ެPͭ8i)/��� �#!�� Jp�"�s�zF�Jݯ�Lܴ�>yl2Gr�j˅b�{0A�c֙�h-�p�T_��]{c��è����T�QDp��4��G�*W�kl��dJ�й�n$2[-�� I ��wI�.p�lK��p�5�0:�t��� :�<�Y'�i�1\�O ���(�Oj�wŇ>�-+s�L5��3*�2yϴ���R#�kw���g�I�oZU�d��;��0�3R?�ePKZ����&�ͥ�HN��l$"_S�dp�L����ӤR�M����B������$pIه��V9�g��Iv��W����?��e�F����w���9����]L[�BUH��F�h6{�/jhH���A`Q��>Dy)�P�yC��Jc��Cv��h�u�N���nFK����d��o�혹����
��xd�$>qZO>�A�?�Q��
u��}C�������\����4��`-C<'�����-��Z#�?많����rx���yr^�dC[S�́o�P�ow/� U�U ��\	�nA�H)/�y�{Q�9�GEj���\D�9Z���7�ܠ��'7?��g-V��,��.a%�J�i��0��H�6������1M��P�#����XH0Ư��]M�0����&�e��E�M�k���HJ��Ѳ_ݰ@L�<f�t�F�_a��U���������'ߎ��*�4�G���Z��|G�X/���:$��KF��O�GT�>�Voƞ
~�i����#+&\d�M�}����!V����S򬘗�-��~Q�t�z��aG�o����;��@3%�<�DX�Cs#@)�h�ۂ��4����O*p�8�p����.�>���{V� hO�	��5��SY)����3I�>:H+-ED}F�I�U?d=n@A��?�*��Y���5t�j�L�=������y�׷��@1�ϋ����C��z���4u���Ճ
:�dY��P���B�5n�╉�M���[�U����&Vcu�"�{��d�!���y�I���辎������Uk��EG �uq[���@������`�~;����'���l7W=�R�����G�rQQ�WhpH�L�ƒT�Z�L��XљU��C�Ju>�o�@�4�@�nX2��.=:�%�Y�t.��8���)��#D}���ro7��\�i��|�B.����/v���󰪦�������P)��fUH�݃��(.�sc�/�*�!�q�m`��HH�z��[&U8̬��1a���[�
1l�"��HdϪ��߼z�v,���iN�]m!g�zWnMܯ9�N]�J��8`�5sw>����]͟��o�^�~����m[�Y��V�=^��q//�*��� ��g�G���>ٔ�}Q�#�EfH�o��:����^ ����0z�aaT,Pl�\�zC:��Zy�.���_�}6�����-��<9������؂��q��I�YQ��+�Ίy���G�ْ�I%x._[8���q�V I&xJ���=��}�Z�ge��+�g�Т����=?���B�,��d;F��Z��t�xm^@�uxfL�������,��܅x����#�����Dz�!V����k"v�΄1ѕ��y��m��R�=^_��|��)�d1dɽ�'�6�����p�˫ar��/�I�����θ:�6��Z���Ȣ�E�a���k�ҟֽ�����8�������P'o"�"i)�m��Aکd�@�V-�5��E�§ա�xV�PI�pB77�����.&�#�B�����v��R[+���c D�^��a}���P��}�"�e,ݍ�/��ё��N��r�i'Z|9�@	���:x寱V��%�yŚL�J�ż�x�EtC�0F5�c���H[άk�/�H�SEx�~��?`��A˂>W/��e�׻y3��$|A�jo �8�X!�@!7~6j���Z�\cX*Y��h�u1F�JB޵Y��0vi�kw�ur�
�j���ȳO0�sb�, ���Y��Z��n������2\���B��,H�M4�9�H@�^3y͔,����D=�~��A3�e21xPD�$ȘMǹ�H��$E�-7��}u�<"�t��Ǽ�%��N^�b @�#���N�)�(�͟���_i��ꗟ���'����+��KMBB\�d7���#9���xAJ�M��%6���F�w(�hQ�M�Cta��e�#�y�"�kq-��%�4��(R>F�|��6�٭]H饭�T������7 �"{�Nr���N�n�n��5 Z��>Y��j�^M�#meX�m�ċX�;�&1�
��4�!��&A^;`\]0��g��jp"c ��&��
�����&���;�C���y^ʻ^�����m�]�|]Xټ-�gj���R,��JW�(`�y�<�ރ��ܺ�V�D���^X����j�K屮`4�(�-�9y�`$�.�i��rӡ
�J¿�#���WhU�fz��Vkù����1���}"�9U�<�J�գ�Hy�g�P�uAJ>*}w�C!��5���y�؋�H�92���ڃi߼�]��ևP������Ê�Oo?��5e��i͂��ϠI����oh�gOi��6P�� �jbgY<���蓔��h����!�9~����d���d+�B�����V��n#`9�C4�N]�z���V0�h��7^��.�}xGQ�[i���x���A�VߟE�FJ�J*�4�����VW%`D�;�>�/��6��ޕco�C�/�Sw�o�ݘf����&�0��<���:Z>H�'��D:���JZА]��ScT&GƓ��}{��^��=������jSh�l�R���\��.��
�k� r|&�h�w��%�a�����jb�C��Z<���#��WO�C[(��1�na���H b��/8L���'��%́�*4�M�z�G$���(�F���N�@M��1C�@��2~!L�<UN��f�S4�׳����f�4����R�4v�,�q�x2�?Ln�>��t�[�Po�-N���6����B����2��[�fJFK�gnPG�o0X�^���Ck�9 kk�,����^o�uH�D���9��ۿY�ij`�	4<Fڱ37ߝ�7y��!C��1��5�����0��G3�'bC��z?�=pw�J�<�j"�["t8�=� ���։�D����G�J��{�B%t�a��X#%u����kжKgF'��ʗ7Zً��]��5K���w�K����.eG�`-9KQ�U=k.	�T�UM�?��{��Q�&�I� �0 z���]S�;����@vp�O��:{VG��p��R,���!3.g��gHY���/�It�ږ����Կ���ZͼJs��HD7���}�0Y,Ɇ�ox�\
YM�� ElO�/%���b���ϙ�S������t�]d�V�u�{f�Ԝ?��@��C��r���:�z�$�/�_.`aI����e���G�/����E{AR#�j�Kz��T�^���'��B��ʸ����Ժ\2Z7FmJ� �o`-f�t:�;QY+��Х�O��]C�cfM��ߖ��WTmz��2;�0Ynh����RM���϶3dĕ�ӎ4�;ݔM�.������A��Փ��}��9�1E���oL�>���L�j�S~}N�~�;z6�/T��qC�4<L��=�x���W�V,>���@@/;s�܌] 34ñB�Ybsm"���E��6�6��g:p���6��K4E)�1udR��e9�9c�GN��.H{���$I݃���<�wVx�~'���{�4�����$�!wGGv[������1�([e�|��B�1��e��������,r�L��!ҕ�y �qF^�:�7K4.���h�jhsi(<���Q���Kߴ�7i��16�[��g��ږ&�1��q��m)x^a�U�x�c�^��.��O��5r�gP��-�}q��%��kO�3�[SS��V4m8Ffw�[M�4���<�m�}�����d:��olYu�qd�,���e�m��~��� ��$�lr�L�g��B��H�?w��iMo�E�Í�q�#
(��'I��'��44jFwéhO$1���E�+�Q����lϊ�O�VdqyP�t�T�*F'S��%d#�ж��M$�}�����H���蚁P��u�O^`j�~)����F� �:���u�	�/����?���@o��t����p���:�|YS*��y� 
۩1��n>�MPnΜb��7c��6�������U��7ΡS�":��*uc�3�Ѯ����Ҕ�oqĩ�401�w�ꆂ�{�����Y�'�o��(h͙��fX�J:ܑD�FM!z��LY��y�^�I���ڔ�W� ̾���N&;���C{��=�~z�����]��*^�����d��[��4��n�&�*��j���lp
��(��ݎ�v.6Ρ��z�GDV��q��{k�ۅﱂC�6���Vx�ME�ߪn��Q�2��buR���˳�1 5m�4�!)�^g��+?y^\n)��-���z�U
L��K�Ǯ^��'�`v�{�u�2��`��|X��F
a�P,�/;��r�*B��<=��:5ځ��Ԕ~X�l��Ԉ�v��3+�M�	��0�1�/6}���I���T`��W�{�°m�0Yc&o~ܑ�D�^P���~B}���[��&X��ZQ�Ji}eV�٬H�æ�w�rF01�M4`/�.�575pH����6��	D�U���1���+�+6���7>�\-_aMz��i��v���4�[e�o����e���'N�����K�]�3�� �"����2�5>b��n8��QD|؅�|���{�~۹T��?6}�c�yP�R-�u��k���ۜ�T ص��r�ǻΤ�@�Xy���^v�o�N�5>�d(��K�uq��ܫ?R��Q7$a7�I����\��9{�~S_�k3���%���<q�-zk}9U���|�ƒ3���\�0��Zz@�X]�ۭQ� ?v�u�-��k����)8^�f�=�Ov"�1X����o۫��Mp@N���R8kw��hH��jD
`���(7��N�W�9L���������>�MAsљ�j��K��L(	�����HH��=y��n���{e������}�`��-����D�D�����U�Q_�W�$i�=���LѠ@�]��	������8fŇ��#�0=b4ar�+��{�*��o�~b�5u[>'4��?X���D{|w�4φ�	���{	�ئX��Hb]��	�{;�b�y�]����y�Q&�̝���x����q�������pF�ݨM�����1Ueʦj�X�Q;[o�z�o�v�އ�
��vr��j�<''(И��N��|�	W}�ŝ	�(�4r�����X�j�'��ΚJ���}o�j3-�W��3�[�G��Rz��etCva��h�Ҏ�>g������Z��\�+(����i�e��B��NE�1�����>�*��L�v�j�#��1a3�sX"���@GKny"�i͊R�W�+ �����n�u�o��-�P%Dm�MJԒ�ċ���"���16�9&wIW��k!C&6��5�,t%��n��J��ڢ*����!�Pɨ}6\�ۦr��j��U��J�ʯ�����#���&-`�V�$�#��:��i@	%\g���￮�R��^@)��A�r��Z���gqQ�� \�������,��D�����$�j�� �L�Tm�c������i��������	�]���O���1.<����v�B�|(J�ȧ!j��V���1}�U�~��8��Ƒn5h��lJ�z@4k4�^%	�i��"C��0��C���Nb�k[fS.�C�С���0ƚ�e�6��Q��eػ�� ���sbu��M4%kr�_��?��\OH�22`N&����@�R�Q�<9,n[_�1䲺93�"1Xc������-�f(sN�[���ĉ�{q��2�q��zr���D������}������H$���O�(�1��k.���N�,��"nm�.�1��K��h}_��֒�i�<�fN���+jԵ�o���q^�9
�-h���)^|*Z��,f���OH	Vtl<<�n-�Q��T�Q'Lط&�?pV�$��$���aۻcQ��eßFE�/�lѾ��i�"��xn�|� ����Zp%�N�l=0�"u:�`��a���m��0�ﳠM��-UV�5%���7�=�F�3�-�Q$��c����Ľ|��ܔ=��K�����n,�D�e�;��~�s���Y������"3Vq�L/�E��l/��x�|���8����v�WܴA)��A}�UZ�����g��2Ș��̥+A]p��5gc'��v7j�X֎��̋v�[�z�?�*�tڅ�g��h�U[X+���iX�����G�:��|�#�|8r�%��>�4F�*��m��/9��	4��<��rM}�Po�����q{B_�@�.�0*��Sr����h�̇�԰������ۂpf�-�<$��_� hkIR+��o���sx�׀F�A������������bZ��1���&Y0A��z!�ى��@NcӾ�ȧ���G�s�D����<�f�Ƙ&$È|�2h�O4�I/6���f�9TE䩍��Z��1�-<þ��<��L�ئf���	��cu�6��A�� ����s�ō&��O��V�3SpVE�WK�3ϒr	�V_��e�\ž��ZPoT��v.4.�s��H�B��6/`j��ފ�aG�A�	{��l����|���f�W[��w��X'�X�r�	`�� �pH�=���C\���K��Y|��%�4�;���ٷsP��3�1�sY�d$���1�7�錜� ,���YՔ?�����	��T�9P���Y�Љ�W�3ꅔ�x�"}q���Luq�p]C����|�����m]!��͂�})��S�K��|U�RX}a$E��`�"��A��N�I��Cz!Za���3	��Ř`�n
E�I���w�n������J[g����C�w�rS�Gz���%�?GtӾuuf�*�$l�|Ç+��F�����3[$�k��)N����%�g|/>��D�.τ�Dp����/�tx]�n���EPD�Mઘ���U�}7��=�+���a�5���Ԥ�e����|T\��������7��N�rr�7�>E:q"��-Q���}�N�n����*��eC�2����K� ����a�<�PK]�f�*j�#���9O�����"���U��~�c}ꌝ�x��zA� �?0�;G2�Q���Zj���-ΫP�M�+�.��@-�߬�	.Q̈��8_a������Ar&7�<�cO�]Q�>���U�p�G+���8#�NH�A&E�V������f�!���%�U���Q��=�C���G�rR�ǽ��1Z�$G~�p��U^�f��J��+���,��/�o�B���T�Y�~�h~
�ò���?��=z�[2��V����'��9�~�T���/��/|=Q�XH�m�%���Gʪ��)�:kv</���@��1P\�,!��X�G#D��ÖVq��۹�[�����b�j�-Mx��}>��e˶���~��)��7�����]B��RQ�kj�`�}f[���2��um&�O����ئ�g���~q8a=ݑG���
�r9Ç��FR���x���[���A���~7Z $�b��H.�r����$�9�Lf�M��D��0=\���'�%�$e����	Θ3sO��oY�iΔ��A��j xJl��8����9�#90$H8� P�1�'4�~"��M��CL��yP��kq�v�'0�	����8�6��_!�f�	d�kCT:�� �>p�M	6�7�;�g25�0�Ӝ�oW���J�d�����ۈ�E�r+�������,
l��Y�������v�Ros����4��o�Ĳ���g9��:�S%���1&�媯\��\f�����LHDǇ�_�O��e�D�zG}k�1ᚼv L�ud�
4�=BM����$u3r�������t�?���>dL9W=��lF�m��{f��m�~JVqҀ��M $���M�$���j�' 49���>g�^��Yh���E�~ P�_ߛm3�m�_���tXL��(�� �ߩ�GZ
4-�(��{,�ǧB��˭�%
��Gg А�j�J\��"�D����Á�_�E�ϵ����z�@�:��A�שid��T�����8d���5�̆2z��VpF�
�x�J� (%Yx*���EDÒR	<Q�V���Փ1�􅿙(Λ�B�U����T�<������6�h�YG3o`C������He�8a���+4������EF�e$1EG�W�jT����'#D�+w8t�?F���l��h�������ٲ�̬mT9�>�h��� �e��_��C�O�'�M�Uɍ�ɏ���NqH�V��5�ˡ�W��m�[�^�*1V�qQM�}�י hۅ-:k�B�=���Lx��-��p��=��Oue�Q�-q�/@��*�Dw�]e?�]���`�=ƺ��.q�e[ #����,��g��\�����z��;>���	D�]�q�҅4͋8�5���9���t,M�:�������g�[��Y��E=�V��QK<Hf�K ��5Z�G����gމ[൚�]p�`��oETG��2�)��s�>�C��r�P�-g��Y�0��ʑ�;�E�B��Qv6��rd�_f�����Y�ԋҏ����~f>i'����>2㙃���!� �2O˪ �����~a�PPCf=�Tx�ږl`^k�b�/�,ƴp��{��l�;����4o�����څ�p�r�~SB`W	@�lf�"�(��X�B.�B��yuh��J�7(��@�]��7���.+�bٸDӴʈu��:U����$��-��8����)�����<�i�v��y�4)��d��'R�4�R�K�"���P��$�>I!OxJ���eX�|Q���70���+�ʇ�s��S�j��x� n��	�O�y�u�	�Y��yn ��X%�����+F�-(�8H���c�R�\�R^D��d���ӴO�pҨ�(\������{@��oV-��eƏ�O�PJ������:���K1��9��0y�m<j���M�a���nq;�����B�x�U�hqu��/i�զ
����k�ԦA(d�s�]�D��^S/��j����g��p	`��=�m����z�Xs:���d���J�y�a��֐ڌ `�P��pvt#���*�?�#C�1��= �*�qu�pm����	#ӗ��?Lm1�L���n�t}>`�()x�%&�q
&(]Q��R�h��l�X����/.� +�����7j��ty�+�]n�4V��=wI�ʞ�:#!N�mt���z��ȝ!y����w�zͽ�y��k�#c�@�.��t��B�=���d�y=���G.c��Ʒ@4�̪b qQ���h;��!�hw;P�Kג娼�Y�F'�2�̴N��}���L O����D��yFD8q��}|HΖi'7J���1�HZ�5�'FD����1����Q�Ժ}I�-���蚬�{e�zK�h�� w$Ԝ|�ʝ�-�s7!&�����
S��1L�e�%������JO6�z�olt��*��Q����"�)1�4�}�cZ�V�N~�N�^���>�W�H5,[׌�o5��
���љ�>� �E};*Z���!z��,���E�;�9J!!S�zN���Phv,g��vp�A!,����.���3`f7�-͔�Ȟ�"ڞ�c���Q�h�!���-����w穕��0C]	��I����J���w�ζ(<n�T��]����r
g�9�y����O�bt�W��G���Ȫܴ��/GĠ]'q~�R�xdT; {��f��W����qy���r���owe1�|<O*%�x
z	8.տ���9
(MVg�Ӧf���YTI�$��P]:��ś�߁�
OL�?���u�ląc9V ��2���^W<E��9�yDF�,�0���E�8v�&���L_� �����յ<��Q{d�P`?=�wyO5�qGl�D���D|�s�)�v9JCG�'��Fw|�.Ҽ������(�Eh#�(HF'E�u1C�A�(F[� &�=R��fYM·�#��q5u�F����k`��;IF��Ѓ?��6(F�}�*g[�jd7���]�`������2޼v��+�Q,����i�������Q�����Ǫ�t��^Y:Fu��|̧Q���ht�`��t��Mh�1��ޓW������?�e%>=z��q������������=���B��:����]�!.�F��TXY�xQ����"Nd ��L�-74=�Ѧ�(��"[�P��o�q��++l[g����I�c*�ܷ��b���m`us�n$@���|;6=�!�6��(��e5�/�Y��+O�wm�$M�I�o (x[8�q		ip�➕bh	����Fy<�̝)\6r��~5ޟ�%�Mo�IF�GK�:���XT���Wq�(�6\�QlV4��6U�@\�Ud�.� ��k��l�R���6�d�	Y7��7S���0���W�����au��U����|)����<�\=BNsr�v�*���� �N�%��@/�Gh��@���%닕�&����W,F��~X��i]<�:u���6������$"�HXA*[(��u	�@z�g ɷ��E9����}C����bp0�Eb�o����g9�[(2��J;�Ųu�K�)��Xn&��]%0�z(bח�/��i!�d�sg��Xc�ep�݄O.��l:�犯k5T��s9�sc�4���nk�낯�t=`ɲ��Gi`�N�F��0���W�N���(�n���� Wl��|�|�g�c�F"�k�������H �\� ��U���z�J�jɜ��?���w��"
�p�o���#�@\�o-�c.������Q�cj G��^���JI��*�Wa����3�ڦ�Ns��ݝ�Ņc��fS����?�D����~�n���A�u����ʾ�a����j���\�<U��h���?�k�{�Nf����ר�ލ�bB7p>m��7f$���a1Ô�r+� ����-1@��P*?�K�<�]#���a�93�?�z��tM	����暏߫IB"{�o���v+�`c�h<m�|���S�R���zj�F%N8��ٷufS��ʣ0�Ȭ�ju"�^
ı�$ ��'�w��{DE�!��_Urn�&'G ��"�����_l"B�b���/�p�O9�Qp��&�w�	�fB��n޺Aub����������m4�(>N]���<G4D�f/� N�'�1��g�4j���suC�K�Y��{�m:aRbs��:�۟'���m���.��F�S���R=�$tИ%� ���0	��u����bu/DZ�-+�
�<ƜEz���nB] �U���xv����+����ʎ[7�&K��¨eb6����A�j(1.�"|�%�9�T���l|���#�rے��2{H�6�/��hmZ���u����'���L�4�����h2�WB��2D�wgMs�3LԖ^�9�X�y��Щ��s�������[Qΰw��[e��v��q�G���	tb&^-���2�����%a|��g���>�`\�4@�v���f�`�Ql~/#�K|�T�(+�S��DiE����IR[�J��cD���8�D1����T��1C����ٴ`��wU�:=�P�O󊂒7�����g�]ܟ�[y(S��
�����(񷮌ڡ��y>�aH����%�U��'�oF�8c<��q�#�G�3wy�����)��x���?׀e�p���Q��2�uA\O�g*Q+��=�sz�{B���R����wBa�������aG�����m�Z�X޳W
��$��-L��w�F�@{&��c-�,�w��z�W��n��/�<4���a-���O={�	�����'q B*K���z�2T�>V�������i>!�GH�G���ȡ{�^ڬ���5XS�V P�1��������Z��J�=�T�}l>P�:)�P�+������Z�J`Tf߲C��KE�6�v�k�Tر�H�>*�X�>
�=b�՛���t�0�h�l0v�۲x������]�&�������o�*"���[�M7Ʊ�����>-����6׌�����|׻�����m�\��ϫ��Y�ubL�`�m�-�,�D�g��0��y~��$�\��&���iɳ� &6=��!l�b�G5�|�z6�f�O�|\���f"WB�c�Ϩk��ʕ�r�\�oW�+�i0s�c)n}�Z�?�[������>�7�@=eHj��4�8�9�9������J����|�<Q���W�1W���{4Q௢A�i�Ϗ����-��9�r'�'���
�;[�,-��$Gꩿ�8/�.ؚ�*s���q�@v�F�83:X
g!��=)��p(ڍCF�A�φ�ֈ�z�td<H%bQ��؜禧OQ0]�~��/]�jv��2f���p�qq^��Ky�|�{��M�->Ќ�Dk��Eks���1�&��� ��Z��.M�C�Kd�����s�������Wq~��v��9n%�HQ�~<L�� ����çX���j'���7Y$Y*����I.d!�x���&d��Bz?w]�͒9���\�/�Q�>�A�*H�&1p�<�NS���V#j�a\[�=�>��|��M�Wn�;؇�?���(� &\6�"���NZ���ާ#t	o�LA�~|�;@g�aK4:�7X�[Ӕ]!���Ⴋ���s��q��s:�b�P��SK���d��0�NfE{�.�'{Tˢ��
 ��~��@pH�=�Π!M�0&]���,����㽵��S�������K�X�?F����e!��ʧ��6_b���q7TvOظ�5�8p7oࣻ�%M&��6�d�����r'�J��?���D>|�9���f�f�; ���t�\��z´$�X����ih6�gޢ�O�3R�X��Ϲ��Q�`w����$�5�=�a��4�rԎ���n����Z��YUmt �V�3y��"���>���
"�tzd��~��(���)pKd��eF/����8.�O�5�FxgDD���)?+U$�pq\��)'4�\����{`������״��s�d�l]�Lx6U3H���O��z���*Qn�E�*��3. �@9���V�[��>��u� ���/���:�\4�¯)�	$P��TG�����B��Ču�#��1�r��W����P��X�t���8����nj���=@`�� 4���H��A'�o���R\��$f	]"1e��(��F�]�0@�1�;)����
Ϧ·�o�PV��Hxn�У��Xƃ.���md�bmh �mgr�ʃ������T6��2s��Md-�ذ�q6CE�]����q�U*��pR�w���B�B�U>qAbDٲ�k�"���|*�{c>�9ڶ�x���Ҥ���8{~��j�l��,�/*�U��3MD9رέz����k
�T���<���o�����o|�t�`��5�?�1�l��� 55�#gؘ��뫂�F��EK{�;3'���%b�Dc2u	��\��RLb/��m��Kf��볣�=�p@4�W�a��a�=嬶!�I���t���W�J�P���fa��I���!b�3|+���_b��Gvp�f���V����7�%?"�֪�G�L�lk�:=�s����Xa�CYL�ydqx8�E�Gz��B[~n�S�|5F|~�E��O�u:��`�f&�1�s;S�����כ�?2���<�����՗$� rY;?�E�����*`�\�u9bvV����~���2	�<Mu���L=H@��2jc��Ek�~쫨������/�P��C�!�>�5�Bџأ����{w v~i.�z�NL�w{��1�W^��Tny����S�g2J)��� �
�秶�y=[?-�#%w�8��)�'Ѿ�Slzi��t��V��W�@^*�4Kn�g����ZV�.B�͈��K݋�Ŭ>�Y��d�d�ش��:�
��m���F�r��8���X��Og�c¼W���z���5,TW8tB��h�� k���'����ۭoZ���i���}c�d�r{��Q�ݎ���q"�0�I�/0���Ep���Ԋ>��1��7�L:���;S�K"}oy�G)T%|T�����iMa�
�~��:�_z���a��zp�(/a�#�e����;eۅ�|�8n����XT�{/2d郪��DK�W*}¥O�$��@�J�_�4��6
���fd���6���ԗӱ�Z�+������!�M(w�"Pst��bی�K
j���*�Y�4'y$V0��lmy��.�w?¶�T�Bs�c�&e��9�EN��E¬��Ka��X4JH ��f�+@�5.;H���dY�a�x�M2w�#y-���&zj1X[��1ͱ�#	8�/��`��;�AZ�o��B�c�i�7�8o���EQN݇���p#w����v�<����攌Kù�7P�̷h6Y	ܨ"ݢ����*��T��x�ߢ��5�C��B��0Nmew�������<pI�]�D�e5�dh�v��n�K�'m�h:��y�����P˗3]U�{e��/D��|�ss�Cp�Z!%ϛbf����n�R��;�����Z%\'�
�fBd5($ƌ�g�X��v��	x���|K���PA$���'.�Hxi��p�R���4��S�5r�.خ���w0�"K�=H��u&Vuhy�ʖ�r�u�m1�(�����w�*7��8|+bݽw,�?=:�3�΢�_
O�z�]k ����*�́f�'P�!	V���:��������Xf�ݸ�7�#n=���f3�17/�����7(1VA2΢�<��H��k�[����#�������t�Zi��-�!٨��BА���6E�w���72%���*�=�n���?��̶
BT_����CP����\1dy��e�@��D�\x��~;��� ̈�ر;WH�s8���	���	�!�k,�v�$$��j���.��FY{":WP��#P�-����d�����$���"�2.o����?�{K+����Tt,�g����,Bv�4#�<?��ʨ�ח[��R��u<Y:p��S���<�_�V���X�#-n�̅5̽3�R�f�Ϸ�f�t.�B�&��(��$�ț^{"�4�!`��Kw����Q�5� s/�?�.Hw��VС8�U>�c���(�)b�3��d�z*Q�菸�œ�5O9e�7���,���vO���L���Zi?σ˜t3m������~�/�Df&��/��嬃�ϫڇ8Q�3R*�=�I<�4��p,��;.������������Cl��2^"Hl��<�E�H���-��U�K�d �Z�����\86L�+atM(X���̮��=^+9v����M�5s7y�_�+�I�E�d�N�vضu,�P7k�οp����5TBw��XB��m
 -1�?��'��#�G�����?V�I�|��ۗ*����y�lk<>џv�ƍ|��h�[_��~,���$bPw�b��N憙q�d�{^#]������!�ߍ]:~����}g"	���=Z)��ʙ:�9���iZx�I~���T�ȹ����B�D�`.U���fr@Bԁ��H��aQL��>[h�?pJaE�a�#HS"�%�m*����t�����mD
auP�=q@�(r7;w.� f��aoSݵ�m�D��M�n���d����C���@�%d`�-�h�']��:�hoSF���z�Ƀ�E
ɯafC|!K��:�p�pH=|���.pB*6����iU�/��+�����Oɖ����x<p�Rv��r7���`�_KjF����E��6��"'O7m�/�2:&�/���T����z6�����B��3�j�jJ7l������|"�3G��V�4�"H��r��L�Rv�����t��1 d�t˞e&��G\�Ijt([�ÝHﰄ�HL�S��C�P@�G;�-J�xCF�̟yz��&�GV#���d�S�����;� ��=��:*��6�����~����#����Or��u.��0ˉ�� Jp֤�IQ@إ�Lu��&���8���7�����4?��W;�@A��".���a���J�z��YA��b�oN%�;���-�Ѧ�2���~3xe�#�A�:�0��������*ӮU&d�u �ţ��Z'.<�������Z�|)�Sc�IC��@U�w.��eb�vZeV�|�s($x�v�lFyg; W��xAҧOL�3 r���6�a����Y�̾�1��?#=Cŀyp�p$N��S�TU��44KM��D�����)G<����	�L����kLY�:Wr�i}*�bOF�Cl���n��Ȍ�3���G�<�ϩ1�"24A��������x��G��q�d��/����:�7���!�g��m2`ljr�[�G��
K]3׈q�¥����i���� � s5���'
�˷�ӎ�������~��*��g�Պ��jO����P!���{�]:M٢'������G#�z���BJ	�߶Ȝ�g(U\�l��vo�����YD��`5��a@�n̄$M�ÇV�-Gi��ak�rN���{}2�c[�m⚁� W�򴊯�q�7�{+»I�)�g���W�e�I�^�2c�1���gRX�����^�V���!�G���*@U9b( I-�n��^I7i�?Q���Ā`mY�By/R-ކ��U�
=xp#F��rv�����j
��kq��v��l�z���h�@)�=�(���vy���T�������1K67�P΢J<3Y�g,Z��� �P���j�AFX)a�Q�f�6T��i�����7�'S� ,n�����Kl�,���%� �2�ZC��T߭^m���;���]����`ԗ�5�Ss��L�J������RV��U�#��94jp���t��ru<ý5�x�չs�㴃�����%( ����������&w�������g�/�U���Ʀ�o{��D����������[�4f��Λ�=�?YL����Wa�
�|��s@j�n*�?f8��C2Iuf0��C�[J��>���}�:�ͻ}#-)��ԭ�1��뿆�'����N��)]���T���S��$�w��~4p�b0I|��kbgM�H�Zrʥ�M�-y�j�b	�/��K�����I����`
Z��1ov��b7�A����	&��5�/F܉B>K��C����������]YjaK{�氷5���H9��m&�H�{;JJ�~���҆I�¯�<���_3�7)�k�Ϊ�J$�����"������ǲ��J,-F���0����ң
��%OIG��HG/�\�{��V�4�ò��(�ML����1���Nz�۔7�l���S�r�sP}Y�T����K �n���Y�S����C��c6[�O�D�P�x��Am���$B��Ed:�a��y������+�xD�Z������)�.󒾣��ּ(�I��"� ���-C��~NTO^�Z�w�#��Bl��v�}��|]V���?Sc?;������C�����W��( �g	p�E��ݭAێn�f���>�7w޷���m3���;���v/�����GѲk
*.w��`�V^������b�.�{��FvB:��3�L��@��hQ�e��.�]��Pl(☐���9䜗y���	f�;�-Ͳnk��Z�A��n2�;OO����$�e�����M���"�T���3Uz��FT@��������b��?ɔ�P���D��kuje|��>�]�t�	�������v�N�&�h�t#m,�n�v�10����pkS�x�u[jf�C�1�������{�2��X7Mx�x&�q"�[u[j��Ti	�0��}�)׼�vm)h�\��x5�E��B�m��<3�ĥY��{������&���$��7�,�1��/Z�hZ��dB���:��C5
8.ӶZ\���F>[���J�\�.��xel�9�=$F`��[Ս�{%�!��PӼG�6�3���^�����Pm�v~�,]�BP�вք�z�����-�K���Э!�����V/kT�����t�`��s�Qt�GK�i%�,��aDA5�I�����,�F�h�U��0�d7dg��^w04�VԸ��l�����u�u�ָ�.��iy�D��w-�g�8�:W��/!�߉�� ��ݨ��l��Ȃ����!������`�,4�'(���lՎ� �T3�'Ha^n���hRV��^��,C�m�+-�u7HĲܢ��^6�7�l�j�d�Z����dw�c �C%i�[ ZR������hĻ���QI���{����r�RtO�Oץ�\��d�l�ş����5���l-k7����,gћ1�w�ٶʄ6�� >� yP�����W�~��()J��9.��	�y���;��)/���P2�B�˰�~���2U���l�Cͦ����t�lRQ�
H#a9��{�x;)u<[�d��J�N�tߘ��q�*��󢁈H�im*���E)��w�W����3���H����?���CE�8X�՘��*�ۻ�vU��'�-#wE��=;�&n� `�5@!M�xp`X��[*��v�r��p
#ykE����*�z}�B��q�&aR���k�9���pv X�}�S^�an ��/��&�;�_�A����|Tx��Ag5�*��q]�ª�<� �e"�Q��9�'�7,��u�wP0���_���GE�Ĩ�m}�5Ut�B�!i�+irYت��lmT�j�A%�����u�L4��疥
���n�#�^a�x��э&��d���t�N��za�i5\Z�ň��l��N~��(22Pb�S���p>��֗�U�a}V�H=q��������)ґ<��E�R{)J�ޑ�7@�P�d)J%>(���k1�$�����K�bK�I�~�UoV�a�#Ļ����8���8'���m`u��h�3�b��F�2F�r{fW�/grM��Yb'{��b��N�⩣-6�ø)["���>���b�"O���� ��P���D���\����z��i�B|dtX��1��`�;(XJ� r>��R�;J���2U��p��V�w���̛EC���eW���Q&��\;�V��$x�.)����C�0��eK-�;8��c1_�A9$��٩m�,jYx7<D�X�F2X�_%�w��l��� TWPW*m��s��`%�m�pB,��I��_
���%��H{�Υ53<���bT�������Crw�1�$��O��i,1��o��1 �u�{�%����\a6m:��)`���<�O�����м%!Va�ٱ)G�M;�|n&7�s�#��|z*;���ܟ�p�ˌ�+2|ÜJ�v�J��5�ˮ�|Յ�oP�40�fM�D1[=I��C�g@ݰrF�c��z�R/�����-��L�P�"�i!NM!��`�@= �}V��Û��w�!q���x`�M���⤠a�S�Q��k�����F�t<8q#�˿���R���o��yg�Yi�E�_5���t@����'�s�o�-%����Bض�h�a�t�5�^��<�O�P2l��!D�5]	�j�/��H�8�);�g dUI�K(����&9%||���}���DG�U(V���T�ӳpWo��PLH��DF �;8�D�<R>�r_"{1y����tg�)8Lf��H�Gf��#�I�Ñ�F�X����]C��p� 1G�Y����ߴ���S��\!����0r��3`���,��P��4|�v�}N��E@�E�ϱ;:�Շ��_�}1Cy������p m����2L0�V��]Hb�G�,ۣ�ǼNN36R_|eRB͐�D�V����ep�K>EB�Еr�U�Ģ�;�|�WP{\��p�� �`����{"� �S���7>�&g��,�qS�=�8��MZ�3�4��J�h=���N|L?kPey�(u"�`����� 2;NV�σ���<ݪ�uS%�֢�{��~�&X����VxD/	}�WO���!�J;���q	f�Tni�̘[3MWd�f/6ȥ	qrd����$D�ty�*�x#�L��<�G ��L. ��]���3_�H���6<�L`�W��n���x	qF���'N���W���긒X쾾����9c���(�2�<J+ʛ|�5BR�GH^a��[^�Y���[uy�9CGJ�8�>��B1jUAXr/���a2y <.����^��_!�qF{���;���Hȵl!�1��N�F>�T;��[BA�!���o����UT25�{�>x
w��1�y�d�)�"[ �S�*n8��O�h�-���m�
04]�y\����t}�w%�L7ߞ/�3�"�����
��u;(j5i��K%�g��9��U�G����9��$�H��ft�n�nY4_8=�T�y:.�q
�0%f�G	�j�7�R��`�s'}.�dL����n���C~Հh���ʚ^0���yFO��*J������(g��k9�$u���ؿH�\i�J��8L \��b$]{��kҩ�e̒�D�p��7�G���T�H3�����b����+�Y�ʯ��:KxD�<dɏJK��h5(�a��C�8�	�Hu�̗�"��k���8⟚��`=|�*�
,@C͊��6�K߼&
��C�71�q¤��x�>�<U�9Ɩ����ϣ�%���b&Do(ܲ�qp������؉��� ���r�ۇ�C%m:�B��P9��ƅ�Z�S��G�>,����?��U@����}!��m��X��])��#�������&�II���H�W���?id|��u�Wֽаf���U�=�&�-���=��R���f�c��վ�|����/�$-�T�8%���������8d��3 �u(��������d�A�1�+Z��
��;'���aÜ�b
���ۯ#Q���w�z3VP��U
F#+��ǒ�$'���A��������#;��|n1�?�Tl�&qC�,fX��t�������P��T���BK������1e��A�`�������$-�+\�<�(1,�I���o�ȠS$��#�Q��}�䌤�0��ȿ=]�o��;h������U��$�^�v�xaFa-���7:�����A�� �i�u*F�e(L��N:Hw�_�Դ�G���F�AF|p�D *O_�my�M�h�mҷ�;�T�cS�Qˁ�����;�&׭ʘ+�#$$_]g�aߧ82������O�"��u�f����{P�l�
Ի����Ҽ[=;�m~4F����M�N��,�Sڦ�gk�c���8ӣ|/�N�^�W/ؠ�@�"㾷�?��Ű7��чD�ۜ��y�c�V`����`���=/�p�3d�mY	��_�I>�r��T��|�7iȶZ[��D���ɠu�MQ��m\�d%�� �v��h���> �~�⺣�L��� )7n֎�k�!h���]N����UC����C̉�jqȍ�+�!`�;�?J��<F���-���k	�����-��2Ij��zf����NZr�5��;��G	C#�Q�y����+���S���k�o��2�"{c�%����ӎ�F<l�Z�F� HA���D����8�Ry�3�/�-a�&�L���A�/d�N�)]�f%�e��F�Ǚ_7-^4c���W��2\����t�;F�������iWT�������wW��Y%�M#ǋ0" ����#U�/�=�a�m�V�W��J���;�N:���_:Cz1ta�/I�(Y����#���=�tSr��^�� ��2��J�?F�Ӂ\Qg��'_���_E(�~��0�h��Q�Z��$�f"�Y���>oP
׺ agy��	G���(�7DǼyf��^[3��G��<kj��������z�&s����&�I֎�Im���B��@�̈9�$��-D�ٖ0�T�e�k�i�
A�*��nW�*x
���\%;�����P?��B�_�k(4L��4�Ͻi#1$����L��l5���)S �e����b2"�S���
��N���éC8�- EJ{��h�no*�VX�.��`�S��'��.���k��bݵe��+�	;x��5�C
i͆y�  �s�m+�C?SS���o8x��v�w�<���˺~k�'��i�^E��>_�Y�/-���)�;8�n���3���^Kð'pؙBf���]C0�X^�+ع�J��X�ɺ��	�%�_l���j�.����"V[����8�ɢr���o�����<�>dl�GN��Io\8vRx��a�ݺ'�wfW����$��T��<9+�f���7^4Y�/�i�g�ʛ���&�pM�����W��kH���c��X�N�i���J���T��N�F���ų�E�gM�6Q�P��)�/��X�+��j�H����Tv������w�4�} ����/����$�4�����ZW�Γ'�]�3��i�fQ��\� ؉��g=2�c�/A8��4�K!��3�����W��~P�QRK�0Ⱥ��usz��r��J�d���?�l3�Kx�S!�������ύhU�;E�����D9c*�H��0#L}�^� �q�WR�,fd�n�gG�Y�GI��ߕ.o.�768,��j!jr��%�+�n�bLΞ��>-�9s呰<��mBx{jJ�WT5
y8?�8�C�>���9���l�¡�Os�Р _ Y���"�2�%�uX�<M���9�� ��-;�=`,Cܸ�+����eVsP�
�1��49�ʤm��D�PJ<��F�E�ɧ^�7̶2ՠ"�-�q&8����v��=��)���~��,�>&�~�M�h�����o�3�	!ob�:�������w=%ʝ�Z$����X�<��Nv�Lߒgˮ	�����Z �ޛ�
zj��6(��^amȘ
��9
7.���Ogk��,����RRUbEVr���r��Ov�?�I�/�e&w�$h��ċ�1���C��$��]�"#���N��'�kN�éz�`YH�#�g,�7�59+B��|���5�=��W,{�u�����lW���<����ы��{��C������}��V-�dK�JۮG>��ק~�+8�y?���]	��1�K�Ҹ��7�>I�nX�7!Ƃ昞,N+Q�^Y�YL�̰~FW*N���c��+,�lRg�_@�<l�"���FW���"b��t�F:V�d�G��2���M�*�J���V����i��^{��΄	HF��B
��ܖz�h#����,�	�e�>޲g�FXn��`�}	���˧׀ftZ*v��z�������ߧ���W�H�t�6B�����L�O-���C�ڣ���k�E�*��� m�/+j� Pd�wZջ������׀�t�K�J,���)�_ؖ���^5:Uv�� ��a���,�Y-8��3�;/�8op��x��$q��Z�i9}�AR15��+���j�r�������>�NG^ʩH0�׈�^�ne�C+d��X2��L~����JA��㉆��-��w���?hg}��0�����T�Hc�4��zw��	�?�R�կ����i'��eȻ�an�\��W�2�2���<�(���.�s��V�=��7f�t�$���;��s��n#$*X�^�ˏ<�O�d���qa��F���H��S���🂰�'�*/��%7��4dG�hEⳈ2K��zʆd4x��,%�_>�K۳F�\��r�V��?j����y�ڛ�t7i>icKu������L���4�"�����L���Ÿn�@@gA����(\�-��qR��i���@U�K���p�
�"�S� T��-�m��d^̯م��i(�/O*��*@�d�mw�Q�p4)���N�C��l@>��;�p��N�EON�n�k㬼�������v�����^��ua��SR$��R�fo�^��Zs���E���!�+睙KղD�ue�'^ln�P�6Ε��'N��g�n��T'Y�'k�_Z+Ղ�efe�)��\IR� m���P�e7����r���$%�&X��^9����h�9��|�[�k9��N�a	Y3��&�/ٷJ��p��y-T�1�|�G�߶��.�<,f�$6DQ�2�m���E�~�|���3C�LpWdٛ��55�0��/A�(�<S[�(�t���_��]�Co���7��w���_^��U�Պ�����o��y�9W�u^�Fe�^���%�nB�+��!`��ve5X���L��$b�IC����|��/�:�k��߱�U%�����\.5ٵ�ex���:�\�*��]�k���x�����c���sE��-E砈�\'�g̳�!2���k[7�#���s�@݆u���'����17u����J i$:z�|����r8�-0�*3���{8���rqy�`-�Xv�:�;8M ҃ٺ���������k'��`娌��dvw�i�X=��ͺ޸W�@�Ť-�֥�t&��a���
'a'��5k)�~n���N�z����Ek�u�ےm��c\6=A/M��j�������6bG�S;Z�p�Q����9q��{�	�� �:!P9Vɰҵs��଀��8�6O;�K{/$pd��V�?f�AfI$*��_V���2ʮ?��}I���?S��	k�������?i�>2x��h3�0���ΰ��D��0��@Y�sKuДF��V��%��{� �@����&N�,s>�jB��M~�ݢ`�± �¼Թ�l�,�+��&��%�~�-�K~gsS{)xYP3{	V����>�8<J����@��8ڎ����	L�p?�\!V>Xv��Q��/2��Ym�)�v� ���U�{�����ه�'	����0�i��9�G��4�Zt��G���H�~�0�e��|���а��Y<�(�r�:jğ�3�`������R��<��!�� F]������A���8ϡO	����3�/��Q��N-�����n
������\�A�����쳅�9:��Rͬ"]-5T�[U��nk,�HS�,;�N�d7CjM1�PƳ��1#U�Ѱ
{�ҋt=�{�刢�`�a��:���z�JΔ�W��?WФFHr%�������|�v)_�Ϊ�\���s
Gr�fN��Y��)䟻��h�W=<0 ���쩋��f0}�:i���w��h�;��'iޡ����.�~�J�L̄�a�$uͥ��~dT��6���9�i'p���ȸ��ߤ�tꗶ}�%j�e������/�f὞��,�*n5�b��+2i(:�锣g���@� dp��*�\����y�3�K�qpL���� ��M��8�u�)�M� advDW�>s�����d�r��7��*"�'|��F�U��FX���s�3����0E�S0/U������i�{�M!A�1c��{o�����w��;���i�a��ű�HZ`ŏ��>���Іc�g�4/O�'p	&��P�0��0�$#�腍�$h��ͶNظzEO����'.�ًbӫD-�v^��h�f��!х�����"�9'�X\C�D��a 3g�|�";u�t�v}/�\���ēpe��ּ3��!�43EQ( ��/8������=�k��D�����9N�9�&U���LBߘ^9L9�a$�����`���s���[L��%$���ѫ�W�~�L+������'
B���X;��շ�\0^��>מ��t����L��3՟+�2u�� ��gSL�^Vl��w�[���Ȋ��j�9�.�zx��/�3�Oz�ϼ��Ա7��q��j�����3tv�;�z�e��$;���@D�ox������q�����|_2��eE��N�SP�)�3܂|�\�����S�+>�!|�s�L�R���|�V���E
��^�L�x�>J�QMN[ms#tA�������?��.�Lt�Ƕ�<� ~a�};�����T1bGP"|[�lu���F|�����1r��4�̑B5����tK<?���G��y�u�W\L��\�W��ݬ��:Y��!�mrw�,ʩ\���$�~�w	p��S�p%��ې�.҈s�R�wdV��S��IwƓ�a�AYF滙���"�.�-uH���!0���(U�]�:�@Į��Y�$U��㕀�ˊ�)R��\�W9�,f��Ogc�b9�K��������`Wilc0���_�]=?�J��4Ƨ�(�P���J3N�����Z���VC���9�=Uj�9�;�X��?��V��F4$t����Ě��I�� �5��cǕ����y�!���F�y���Cy�OI�����&e�P���2"��=�w�N�bb1s=n��,��E����l�^ɂ�z՜����|��=1��h��;T]��I�8�%��.
�"�i�~�Hڻ]Rbв���[ʧ�5��w���x7j<~�߫]ΩI3�.r�~:���ӊ� ��+v)�%������'����M��X�8n'�7~'x;��[�DD���w�)��de�v����gX�?�&�c���m��8;��5���G7���ڕ@����;\���Vȍ���(�~��(��č!��s���tb�NQq���5S?��N�q��E��F,��٘k�H�(WE�R����o�'�i'�s�%:�0i���ަx��k��<��# �_Q��P:*���J٬� ����[���N���7~�E���yD�����<e�*�Qc��e�d�Ǝ�P)�Fxڤ��8�e���s��v\Q�o;�b���ċ��SՈ�dU�Hn��ܾ�qX���%�
g���ىcԜJi	��P���sA�!�Q��:����J�|`��
a1ż�����
<ת���Ӌ�U�@����> 9ZI�X��w��S��;��2sc9�_�����vaʠXg�zɓ�4�V5������0�ȯ,��L�闁�߉�$�A���Qh�����(C��P$̺�Bp�UBؔ�ƈ|1� ��T�l��=�����F�X��V�qV�^4�=���QF����|A:bq��8s��e��*#.���x��,�ר\}`������g}����@����:\a����ƕ
S�(Wr3\K�$���4������ve�V�:��|����Z�K���q��G�Ys�d�|�8����m�"�����|�Ita��ȃKr/I�ë�Ka��7|��J��g�,���+Wΰ�,T�-�����D�L)�_.##��;)���22���TE�!���g%�$�{x��c�s������[,�LoBBcB�h�G�.�-E*�����e�=�p���ަ�/抪a���&�7�B��s��:��z���P�Ψ󰵥����QE{�@������ lRTƣ|ȃ��w�|����p���ׂB�1�Fw� N.0>3cA?EGд�)��.u�v쓀-Ҙ�@�ٴ�c�7jx��O�c��*U��
��<�C<�ڕ�$ۺ���[��"�U+ԡ�A�2�֮RǬ|(���lDy��O�jVCP�-8>�IY�Hf���C�&����G�$���"�D�M���v6Dq2(:�K�u��3A"s7�iS�Y��~�q��mv�d��|X�r����c�4��-��<�(V��p�����N~�řІU�i�3��$ݬ�F�::�|R��Q�ʷ'�7����Q%/,c�D�-��
_H�&��*���X�:�,����U�K�r��P�W�������St��Q��JA*����w��J��%_�v.D�Ia[���vy�o�H~����9OJv����ҠW�P#�'#<�ʢ�bG��i$�k��`*��)0��e=���b5C4�l�P@�|LD�+ËE5#�O����>|H�Tt<^^0;��i���]����Q�yp�� �S>�hZ��.�p�8���84tik�ܬ�{��W�m�!���9�N�k�+�GE���\��ޏ�Gu�F����ű� ���~�ZM�}��\!:�y��9�{�]�dV���(�
C��Mqw��e ����wv��<�P����}���F�s�3{�^�c�;��uyi�̎>r�\ đ`!�Xۛ߫ä��=A��t4F��q1���P���U��A���O�u]��j���n:'ߡ�n_��K�@�� .�^T(�:��z���rce�O-��7����^YȢ۬L���z+�E��ԟ;�;��A�+�#���}�(_[#��D�!6���?�l�YT�x' *O��k�Oh��U�O��01���.���6�I�Ou2��Y��[�--��"@����c����L`'45(�r��� �;�&TC?Y}D���G	3�"�.��5��cJ��UIణ{����d{�v(,�kԡ�s�m`�s8ܦXG���r���� fO��]��,RC�>nF/��!�����8�qt��K�az����P��4��bSĸ���n	臭{��^�1��?��'e��;׺���Zӽ����U�Ȑ��&����-�c�UD���X����0٥Yp���\�u��]u�|���Q+���~Q9���)����(�;Rb%��(��n�GY���z�ϗ�U�\����o�2Rh0(ڡf�?7�&|W���
�&e>�ٟ�
�����!&���"&���4�����fmR�O_�0	<g@
&)w6��\�S��&�hAfT����;�/]���}d����'�΍�~uh0m�y�F���o�3�G�f!�_��H���j!��굡՜2�:
�-���M�,B:����	7*K���`EQ-[S+�\/�=����&��2V�o�yLO%y�� M-ڰк�����>�[�p'�%Q׼�� E��G�{7"@��"��4Dh�����8���a�Ӑ݋7cc�;�f��Q�DD>AJ���d!�ebA�Ǘe��WQ��+��#)-�2��m��C�
S��óT���~5u>�C�	�X�P����`5���X|�nt�ҧy���Y<_���rS�T����i��m���������E�DR�M�(��R㍟�E�OU¿�ܤ���Q{�Yr�B��{$o=���!���������h��j���3N@��O{^
붿����r�d� ���yAF�,�i�V,F�����d�NS��YM�#�zSg������i����-��J�|�'�
w����1夔�(:�R� ��h����YP<��T�A����̳�i����'�V��AP����Qb�T�m��$�d=�%�\�Lv����:����Ȗ�Dd�w\.�u6>���'�JFD�E�zVvA�-��}ELA�Z��R�3Tōz� ��2�����S}�@D�o�A��h?o�9L��&�%8"5N{�}+�b��nx:	q��'P)y��Ld�ъ�V��G���w�!��F3��uP�_�f:�����?��P4$a}��p��#6���1�����::z���"F�$��_K8%�~U+Q�n#&|��B�Z%.������P%A�T�8��[Z���*��lH���,�y���. ���Uf��+�t]���q�>a�,A�x����֩Ra�&��A�F��:J�~���o�w���������PeA���y��>�A�W�"4�\���y�';:���$�wo����n
������~��DQ�$��#��Ƽ(я	�=�Ի\f*ϊ��@���km�-�57���_�O���Gc��Ó���]x���QQH�-�ʚ�M<��G�T�Qz<O�n�5�8��l邧��� Ì���1��<	��7TUʵ{r���9��CpgI@�"'	�����e>1���x��<��m}��z��ϱP_�	�3W�l@�7�26�1��?_�1F*�`�;�5�����d�W-���s��uI�к'%�����r����*�"��G�շ������C���Cx���`�2{�L�+�*�D�4���7ޭ�ig�b���}��%j�Ѥ<�Ӈ�2W���yj��%����#������
���}'�nG1�-@iٮ(O���_���2f�>R�X6������"z^�?��fM�#-����)鏿�Z `�p!���ڰo����4��I��?��=� �>n�Bpx(yꛕ��jfݿ��������F�����E���1_����ٸE>y�;�(f��BGp��X��)���5�I�6��_qǂ������Z�Ga��#ݩ������0L>������w�Cde��#��Iyf�=cuF�w�"��p��=��������C��˯�d��Wm��	r����ч��G��B,=1*�ؿJ&�h��0ª��.�`�,3"��*�ȝ�=({������ڪ��*�4��w�@�3���w!
��?�H𦞐�.C���λ��"�����2z�rg���y��「+��E���DA�<u��c�g#�.�ċ��k$Δ�;4��c\můbe���ĝ	�H�Eˍ~�lۜy}�G���1�`�����贯ةa'r�eg�r�Ӥ����>�}�w�(�ST��4�h��[�2��%u��D�ȩ�;0ɊH��x�֩����X��eJ)y�㎷��
刹����+��Z����D(�9S��_�����9���;�6�4�C6C=�O�0%Z�I8*c����.x\"'Y-j}�9^�8ΐ7���	)�1�W~��I?G�������A��6�X�0��`r�E\�v��6�M>%O,A[���}1bw��/\HE<�p�k�����K�H�ߵ�r���6m���J��;��Up�9���P�Q�Rę>L#|�7�w�3;,R=�NŠo��I4	���I�B���H�w���' V�'#��UrY�ٴ����+�u�g9�";JF�Fn_�Q[q�-�D��,/��T��-��"H�D} ��n�����3�y�c����Dm9���.�I�����R^�]:��T�Xǆ�ɉw2ti�]�P��V�cعi��A�eO���҆��B�B�v�'����Q�{��[<$��%D�;�c%FnZ�9���q�+	qD�ެO�K�Fhk�}u~�p�*�|��.�y��8U�^,V�"�3_y���9M7��J���ԗZ�&Q��r�0�g�6�Q)-F�{��� m����o�w��Ť���
;��t|�ͦn���{��Ȧ�/�旚t+l��8�f�R�V��4Ֆ��s��/ۍS)¯;�Nd?���"?��K�
�*�L-��U�f���2��w�JM��+�9�(^s~oR�8�|͖d��R
�R��1��Q~`������خba�����D"4�ց����7)�H�2muj�y�]~+zX�=�Q���@�]��߲�A�&н;�힇G���9<��Via�������t3�eJ�BN�Lɼ��S؉s�l�X������h��F�8_�,���Ǹ�����fA��R{ـ쓟��|�}��a���1*����~wb�p5�3���{���>.F~>�F�w�@U�(G��r��9�T��ˑ�sw�Ba��~jSZ�& &b["� �)��ŎȀ�K��ہfz�8��;�y��0J���7�ٽ �4G!�9A����H��`!ת�N4���w��Pi%}�c���@��d�I�	zeJ/ˠ�j�!��><@��0�]�0|n�K��� Q�ާ%� �UUv����e��6,U+�����
|�'p�������,�ɼ��SCM`�L� 0�I}k)�M+xO���!@-6L	����)�y����# Û�5O�;�����{�+R�R�g�`�M,e�ۋ��f�����p߁<%�4da��ˎ�bQ�>��B��T���?�j�ˋ�2È҄��mu6�pQ0{#ؙ�r��#�a5�F�2�S�kH�������X� .���Z��WK����8�Z��)����`H��CZId�u��_�F�"/
�E<��Ӣ�#��#����f�o%K ^٘ʙV���R"T�c�{LL�@�zdE�n�J��P��J�]r18�[��p?DX�Z&Գ/U������&�b�4xm����,��\E�	O��^췿
qB��x�)���8]\ޢ�[�_��˔Ԥ���߁c��6z�;jA=��ǤI
B:4o|+��q(r���ʚ��3O�����Nou��T��#U$��K\�d�K��h�R��^g9-�J��eE]_��/ry?��Asbm�'���,��v��u$x�q��v\�~2�E�����	6[�N&��d�͑|�$~Ϣp_J{t���ܝT$Nm%$w֒_����;)�\�v��HQ7�_#kV�21��w����Ay�Hz�H�o=`hs�9̅�F4w�N�G*�12�����EA�	i��D��(���b8��j�ÒN�i�!#7��ē�TPEuBU{�w-Y�5:��T��>�АŖE�Y��O�	��%���;�_J��_Y[?]��?O���G=dv�UFY�U,5c� �َ?�θ��n��w��^���9�u�߇n�!��������J������r���(�ܹ@��.�V�Sp�}cT�H��([��������w��S�ol���I��o�K���9TY ���ד���Xb]�s��E���Tr1@�[�-ᾳ�U?,��2��U-�cK�9��ˑ��^l�v��}7���5 �p��<��Ԭ#���j֜C�c����N:1Z	K���_H�,�Sz0�ø��@��������vG�g��v������N>��'�P(Ԩ|�3��Y�Ûw�o6+Gt0�e�ƣ
dN#C���� �kT�usٮ]�'����N=�����Z5	�H/h�����#���Ľ��.�g�Y�5V�NR4�^�Ƒ��mN_QG�4֡�'.��{Dע�G�j�&i���r��9����)h��S!�P��뾏����Z��4�����a�?�j�R�����q���
*b��Z��.�a�sa8���+¨������1�K��S�~�>&9��)E�Hz��+�YȔ��F��/��x��\(W�W��,�ա��4�!z�[Ԩ��}]K��	�ּ�zfگ(vzK��\9�����$>C����MZ��TV�^r�|�*f���>[�I?/z#��~1�֋��ҧ%����S�Or�X��N�ᤫ`����3ȫ��}+�<�r����Gv��V�m�F�`�z�����C
3��&Ѐ�l*�[x ����ޙ�x�b	����ɏ C�
�5���q'ȉ|4:eFm�3�Qw
z@��؂��m�6hΰ�9_̡`V����˚O�ǵ�VWNZš}�� �������"����7zG��1��'n3���#�g�[�4`=��`���jF7��3K&|��Vȏ\ǽ�\�K�r��\w`��t(8=;gˏM�x
���6F���:4|�rW�TS|�]PL-[��R�\�� '6�D�0w-�\��z!	Ve(��͗�*��� ?�$���A�����0�������bx���Z��`0��>H��^FC��D0���V�+�+�IY�)�y�uzu�A 1�`��*�)@���rz�m�N[U3�^��=�MJ=�k��7�W��H��Q7�����B�v�߼.�6�L�z�mۼ9�(fU�����.B�k�����D:K}5h�J�+R�p��"�%H�� ��֬�)pO��A�zj��w���cgP�)?bJ�Ў^��T>��GP!p�p��2���tn���i��X�3P�ݑm����dBBn�4��J��m�!�U^&rYB@Ӯn&ǴN5~��<��l��;"A���*�y�K�ʑ7����Dܤ1���.j�z�;�I���eR����4���Q@ILM��35�L�L���!3?<A��=m���Y��LZ��Q/�fO��OYZ�=��c�W|)�;!��������d�Cx(&7�L�{���"p}�W$Q4������KxW��7pa�X�(hҖ�����~��	�,ۭYH����ǈ�����~W�H�@?���+��}8Y�踻����.}~�0'f�_V��3���+R�*����6��,/uh���*����7P�qY�+�d��to$J� =�eK�I��F��h�ј�"�I��B�1B<:֢���{;�rE�/��Qk'��q��h2������?Յ3x��@�_����m:uK��/D%;�׷�4j#�/�a߹�;}�����ShÝ[o�{��=�v�j )�դJ�Ԏ�B߈쏉��İ��|%�;�?�Y��&�C(}�kPC�wӠ!�
�+��s�W���i4r���m���m�lF�*�bLV�ģ��*��{��)�XT�^���D�*N-/��a>��������C�'�i�I���ʋ��]��|�����Nv�"PgW��������A���$t�G���F���rx���Y_)��f��m��/a��G�mZVz�
L%�mܿ7�+'���r����a4E����Ͼ�����bn����o�)��H�4���v#Ptf���]��$��p3)�{�y��%�T�l�mc���<�EE-G�z�\�\3Ս�����oV�i�Ч��/n�Z��͒�kSԕ�y:�M��U�N���d6!��o� 4�筡0d��pU�L4��Z�9�qAT����_�{�����\1=a�0�%EcC�n�?L��C!�(Tc'D��j��-���(�/d��� ��>�0,�<��h�*�@z�=a����$�o�J���~U|�/����DX:��M����N�Gl�����cw���o��T�ذU�]Gv�r"��Q�6V$�37(��d�uVdM��[���S�^$ع�
�\��m3t�9[�7�X�v�=<��k⡹-M�\e7Oq5e��e���M& �z,���'�ڦ�Q-�M�c�+�4�6�<�Ξ�W��T���뢧caʐ� EI5��ܶ�KYw�l���=EuBEb{~�Ok�˭�{<��*u��D?�Ct��-|O��T
<() f���X�fp�����2�3���|��ar'�}
�;bJ�����<���Q$�L�+���6o�N�/��2-�6$�!�$8?�4��/�w�=BX�Pº#�Wb>�J�Z�L6��J�ޓ�(�q��S�Rh�d�u��[%w���(�����^xf�h�$��2��7�f�����J`�#;�󭞅u�*��︐1d�\������K6��t����of���ox��#R��Zc�[t�K�3��&Ƃ����A~�K���K��!�̿˅�`T4=�qoPB��8"�SC���f�z�7>茺�ʡ���[l�?�'^��|&��}B�V�)�n���,q�ߙ:��쁳����b�4�5~u����5;���{�Q)ߣ՟/���c@�F���P9�W�mK/���8�K���LP8���-JwN��_h$�>����k��C�b�y{�y�;_y� �^y#�婏Y��c�N����>�կ'b�x]��
�'%X.J:� �8�	G7����4�&/���
8�%Ê+��y��$��d٠_n{�@��E���6�ú|��B�0Yc\s��3L\ ��X(p��s1/��
j���7Ɂ_�kb���I䋢z֞u��@W&Fs^}Hh��i� �)ݣ�Bw�YZ�WQ� @ҬÓz��������7u�^�����X���':�m3��Zm�P_d�- G2u�(���(f�ߪ&�Grĺ���Y��K��-��Λo<`8R�S)N��BE"��"����ٱu8�a,\�C\k�ݹN`�?�}w$����rֳ�����`�C�w2����[8��6L~�K�0^��ƻ�n ��������F� Q�Z��	<�e߶�i�=��� �a��
��-<Wo#���YL��]cN��<��z3�_�*�Jy��	$�Թ��io&��Ĭi",�ϛ�<��{6'!{����kZ��3#�g�8��7%��_�����o�n�����x�A�wi���'�aN���x�,�릕����Z�9���:�I� ���$B�ġ?�l�O��i��Z^xݰ�f�}nq(R#�=T3���[��+��U���/�~��W�����n�$F������YK��3q\�.ᖍ�{�Zkz}���T����C����;���t磨ѽ�n�F1ɓ��O>z;���]*�q�塯����v��s�����5��eT~�A+S
�VĎ��e���X������=a�n(}i�⎱-Lp6m}���<���Tk�H� ��ӓwZ��V��%���R�J�q��^�r*q�'|]&���ε�U:��:�������Ɣ������V�	 ��|��\��
 =�1�y�*�A/���T^�(�nz!�J�'�[�3Z_���A�QN�-�*�E�#K-�t}f���6PuT]PA�L4d5��*���U@���`pm1L��1c���'K@ɱ`��*<7'��I��3Xo�ݖ�$/'���؍�)���ʻ��|e3n�=�g���l3��g{����0	������)��'u������X����@�v�h�W�ن�P�a��[8;�#⺛��J�D1É���'�b� ԆF��[�5�����w���K���ËM��C��5L�3�W�;���C�smgV
&�����@M�Ac��!��#����%����aP&���`�y�������8����n�K�(s���|$���*v1
>�}�[��^^L0���l��a&>�'�Giz�J{<N_�A�4m�8�9�j��7�h�F����Pb�����@�����_����ֶ~-=.J��W	E��0����<����>7b�_��5e�8g�-���D�ED���Șll�{X���g<�)W5Ʈ��_���%
m� ��8q�u|���`a<O��*.2��U�<J��|wB����K�* B��kb�0�2꼫cc�QB�5#YzZt�U�-t�B@y��6����^	�� �ΐ��L�	E��n�zH��y���;�t��as'�xĿn
{���ݾՈ�o��3\�5~��dZw�H��C��Pd��z\�U!хb��-T��1<�RG�1���iBQ�g�w���e��gn
X�KJ��(���3l8��S?,�F�0���t.�gL� �c�v�	���r�����B��"�E��� ���~��i�;��Rʺ{i��Ì\F������I#v������ǼtN���K�Q�k���o:h��H���P��f+Ih�gc���ȉs"s[�M�8 �O�-�w@�Oѯz@�����4�Ne$�Ѽ�P��}�}<t�ܸʑ ���j�S� PO����(=@��?#m�>�a Ħ��}��m>}�1��OA�BT��͹��ߺ�8���~�h�W�ʦ$Ƥ�'��@����ɟ�7�jU���^������("� +fr�k�YO�#�������y�&}��\\�Po��ܺ�3-���F��;�V�ӵlBb����Ma��њ�t/�ߧ��^��Q��u���X�b\��NVd���34
,`��,Ɛ�Z�W���	G}3G�p.x��5���[���������.���f��z�OJp/�9����3���G������x�m�f�c�3{-�P!1-�2l˝I|�kl�������bt��G�i��~��u�*8a��N�5�(�� �����׆�:��K���t����*�" A���!�O�(]�V�q��ˇv��{��גQ?�Ç#3%#���-X��7�leXy�E��i!�:��!��,�K%}T��k��~�襆��V}� ��!O+ր��ߑ$f���+8 �s��u��v�������5{���m�7�n�$��,��X���s�DD��_�J}��_�i;Ƣ������g���ɖ�ǝZ'Q�Gا�=<V�˫�2_���Lo����i�u����N�c:�L\���={M,%�}�f)m���]Dc/:� ���j�K�>KZIb�!p��({���̆�� ������60��n�j���#�m���d�&b�Vz`Y�-�m�,'��\�r�=;�T�O�)��=#�cit�9blvtSȿB��_�sw,�+��������Cܱ>�o�7�R�I���ρU���Ozҕ��%��V���iL+������`���a���˵2�D^�m|c�mj����sq�����8ut���H��|�����%�~S��8 )��T�֮M�N�T�����i���."�o1D��������ؾufF	N�R:Q�;ܒ��(_H81��Z���b��λ��4�Ѻ�wM/�~ڢɷ�Pp�y�Z�nY�[�,P�2M���(��!���Ր�1X��VU|�G.�?�{���W�G�m|���sM�w䇄'͘P=�� �B
��j���G^Yo��#�]V��O��]�Y�ްZ�C�M(���FD���/n��o�n?���z$ R����N��v\���E2��eL�H)j��;���a�j��0`P[��Ck���%	���v �h�vH�G�A?Tm7����}f3��.���`���>�Q�79�.��=��9Վ�E�܍���mL`^8_�V�W�(�i�-6�l�0l�╃�t��`�.T������;��!��"��#��z������Pb_��;��pH믬�n�7���j��'���Z��/�.���!�R���@4�
��
F�h�S[����0(9(k�����_@`�]�YL�4�C5Т]�I�6����{h�y�_��� ϰ���r|$�65W�����x.�O��S��C��q^	f�T�=ӛ�X����]��\���.��=��d�Wɽ��:zYC �l���0��oA����fiq���������
�G��³�w�U8���_@��#`i�p8g�מ��<�����³�lU�&L�)��OtW�mC i"gnH<
'l,��`��""�R��I%��mCy���BY��)G�;�"-F�I3M��Ǆ�#Y�BT��
�:�?�q��6�ֳ��F���W�;!dLyxg�[��"�N�MJ�dT��D��ܹЭ��ƶ`�����~�3�$h�^�OT֤[����X"�{���v?�����]ë�Xy��-K�b7��:[�wɵd�a����wx(��/��/��;s'�"�����9�x# ѧq���`�WA����N�H�Av����g�����K�I�θ�E����Y6+z�WfI�fH��4�<�12��Q�Ѫx/jL8P���13�N�ހ��G䣕����:��N�AV�)��YBZ�&���mg^/mG�����0��Co~j�t_������q:��
C�86<:M!�jk;7�Ȧ���mupn-P��;�P��[v������o#���%�vqnAd|��`Zw�c mW�gm�ha.J�5B!!���ʵ�q~�޹�b䍈T����+�d�" ���K{{o�U?��,������c/�<3c��b��)�p;�/z�t\W�����i]��?����8�#��V�Ȭ�TsN�{D�:�7F8V�'�h~f"+E��LFEP�M��1+)��H|#.�,��$�2O:�����ӧQ���q���y
�	�5��^C{�L ��t�4v�����Wh���f:�5c~^-W��#���5��ߤJ����[���"!
���
ط��4���C�U��R��=��
�;�ՊN���i�.�S�o��{�o��I?+�mTR�WW�5�9��Î�ܶ��r�|�*T�I�X]0��Ymv�s���!�?DvV�jx���N����2�ߕ(X��d��畀Y�i��~�g@CƝ� �O���|�]b�tB���:�bW��'6�Zk��%3�)������o]Y���5��\����ZnFU�C���nK��Y�d�O ~e�R'y�(h�H�4Z�gd�JV����ۮ��#���T&�[!�i3�jZ�W�eK@���u/�udM����e�Ks���h��gFR6>8�A9��>N������H�p����UUI�Ԓ�+<_�zT|��F��"�`L���]���:�;=�w�ޔ��5��˂�\
deBC߁��׵�g���$��-�|��J��]>��Q�c>OUPD����~��FV����8�w�v�̻U"B�v%c�BM��E<�IiE�������rg�/k��`�0ń�/lU����˦��lD8'4�醌X=�w�;��]��F�nw ������J*_Z�R�Uut3YA�ZU��HMg	`�i���޳; �������K�������G�2���p�B-t�lo�n긋P�cH8�_"Q����3�,d����CBڅ��8����E�J�U�.�o~���Ɓg�����[��+~(cn,�	y%Z��A�����<���I����zɉ��A�
N���.��TuD}�W�J�����{�j�2Q~��Ra>��f،`l��Z��m�Za�s�г��o�Ck���tyh��ck��⎚t�z�1����B��N�.3�0yK���}D��j!����}�6�Ԅ�ۺ������������V�?ů�k�X7��smXD��EP�z�^i!�c��m�(enK��C����r���^RJZ��$W�<#s��#�64:͇i��� 8j��>白�']�o����Y�8ri��d����|�Y�wj��0�~LЎ���D�<-�`����k��7�	l����C��T��b�d�N/m�������Y�a���}K��Ҟ,�j{���l��5�������_���N��XK��~u��`�Qi������bNn�z8<����ɲ�vvF�W�4��Nuy��5&:������P)@��CJ��E~P�kl�F0���.�6����I����v5����3Ԙ,J�ar�Ia"$����>���Zk>��#���q�p��@'ͨT�b�����@w=���t�f6�l�z�?�r^0�D�ٽ�~���M���r5��+��x�M�F���]�^�H~|�|Cca���0��:m�o�.��zBm]�aT�e�,Qk�?�(A��/ȼb����=�F�m�h ���2�>C���|R#;,9�����Eצ%�둴r�e�Q�ǁou�8�2�r�>�O+����S�����|�x�~�h����A&
u���,��S����U�tj5�o��9�yO�:g9F����4K
l�+�o;O��r�� ڐ'��Q-������2Vv-�W|�UG-տ7]������q�Z��dbst�4�ǘ���}V�\�ctj��I}yr�� >���s@�_wbkm�h)�7�d���{��=�R�*t,�c������4b��7��~e��iiF��q�r�c�D2� �z)��� _U}^_�����8@MYŮ�g£D ��EAm�w��HA�����&.�v�'4�Z�>dp/�a����=���s��*[�o5\�mm�yph"F�cA��%ծ�$�}&���?돷*"��jt8zp�O��*\����{�6�y�X���EWm���吶���d�CYU��>Y�aH�������mjkT[��-�!��1T  ���*�i��zy����S�E˄�ߘ!11������`H7����@��핪�ئ���W%�)���Z��M衭Y��`���m�%$;�Al�,��e�c�?��X���,��Rj�'�
j��K'�����>��aby�䀘/�L"�.ޞ�Lkr,�� �z�C$�d�N�Ţ4� �i�8&	ꄕC���3=;�;(�dUD�Ƣ!��ָ	�75.Y4��:N��ڕ�����ۨ+�i^�؀X>�N��
�������ǡu�gF|#G�(lXۘ�;� ��)��6=�����*X�=��r:^Yv�!ŉ�F,x������r]�h�"�1��@�~�N0Lכ���C�<��	�������5�zՑ���2+9���4gr��F�2r��r�-#�a;xl�9L�l�.a�D�0G_HUq򼪷� �ǿQ�[��$V��_��b���~�b�'�gvC�_����3дz�;yO��f�o�B����J��#���p�����OKd,�����*|C�`�H��)Tq���?:?��P�1��Ћo����w0P�n JLh�F���Ec�9,V�1��`���S�~���҂���:W*���L!�T���$Ɂ�SVb���H Bd���H?PIO��p�ÙDI��g�_�͵�>�v�xZ�vb���B��s�U+�����5^SU��\����y��j�n�c�WS^�FV}����!�;˩Fdgz��{}�0Kq�,.�1�D.6r|>1r�Y3)>�t��y����_�����w��Uj�d��mQ���𝌮���8F��Q��(���x�9L'>/_\4{�^��o�C�O��"$(`����MS0.=y}�MMG�5�~��3�cK �����a�s��e��I���
&�"�������YI���l��TXҩ����3�v&%�H���i>��l�x>�_����vd��J��6���4Ycvr_|4Ys���9������o�[,��.�$�i
�[�D�[��Q���)�z���Ҵ�k,��%7�.��̣{�e�֛u����_�d[S�'��ck]^�J�y:�L޳�	t�K��(��o����?zl�V2����Tr�A�~�DF�6��2�]�B��#C�`�/�"\�胆1�k2,��NH��o��P���M��h/�r]�K�i��S9���{�dAnG[c}
�v�r���$�63u�i@�ëjĳ��B��06��d����Qjy�3O���r�w�[ek� ��8�����f�`ns(�\%˹�M�?U��9�h��WW�������q��,y3v0S�W�l�ˡ�&���eO���d�ԄM"�������m^׮!�����νγ	Ji�M�I��5�!���enH�@�@9D0�]N��#��0#..��k�yvP;(+�5�:Н�D�@��ݪa�#|�a���y��Z�=�<�����%�y���B>\y7�E�L�G��[Y�S�$��`��|�[���>C�5Jen>���O��aҊ��
 2�P� ���\W<1Z>v� *H���e`�B��u��"q"TD�c��"]@1Չ�"��ʞ��n��T �w�w��-�N�o�V{E%�4��Y�غq�UOΎ����L>ˏm杣���o\���z���A���,�r
޺;x���dן|�����Z�Yp��6�D���^Z�����<�|02�=�Nt�I���)�#F�p]Fr��-7(����`~A�c����oB��u��5R���e��1Y3�u�
�AR�m�2�r��|1_�۔�j�r��vj�%Rq�۟�ͅ�Zl։�:o�pt��2�0�Z���U��eiI_�K����'gBP�8m�;�D�պ�Qp�W��qF�B�(o{����1�"{�Rop��ڱ��dI�����׽�e_�xF�WJ_�.p��P���[�(!s)��S�nF ��7a�(1�8x�lU�S��-��Թ�DH��Ǆ�]VX)����-NA�!��<���8��[A�����v������Ť�_�t������a���"ʤ�xՃ�FY� �~��6v�]W����m�h�a9�ba�ΓՄ1ҞǢ��!i_D��O�Qz��H�~��/(������j�h�eFD��8%<�f��g]����pWd{�Fh�7���|4<L�K8H�����7'�a�4��d�J�B�ޫN�rN�γ�%R��������3J�x�u�6�Vz^c�*����_&[��X�a�7>C��޻
�9�xՌ9�%W�u8��ѝu�]�<& �l%U�d]X�=\���5�x��g�U4~`q|IN��wdr�0���|��d���&|o46
2����HsBm/�y�U�F���Y�u�S����W{E��9,S��*3�[)	������R����Qk�o��Ǐx,�����A��N������2=`Iz�~�Lܥc^���@y.F��}6��Ӝ�ߣc@��^�IY_o�a�����N��z��{��r���H�7��/�GG�¤m�T��ޕ���=��U���=䱪����@�G1dHJ��v�0_��j��(t��-�;Hl@�e������1�=��w�(�[ƅ�K;O(&��!�{> �����t�8���BI��,ESw�m�K��$���?���x������� A+>B��`]��r/%�*yj
��76�����,u��Rd���u�������4��aS�r��q�3��~ʘA�nm�=� �SY�����o�du��=[���Yn�`��u�L6S{x�7��{a�ɶ����I[d�k����yn�5ɚg��{�i����l��i�;�ox�˵��G;{����+�)�o��|&)�#��༤��Ut60�G �C8�9y���7�m0<c�K�Τ?�:�ٿ5�S	��Mh��{U�g ���xh&�z�E%~�v߇�ܶ�(?@�0r��F�L�?�L�ڗ�T���,���~�����B`p�JB=�-�8�w�> ˶g��o��<�"`����|.M����
�Xl�^Az��3���'���e�'t��V.{7!�j �>V(k]<�%��� (� "l�b8t�_��F�0��n����}>�w�A��I�����N���%�t>+��@HZ��P��Mm�����wV@�� ���X�Lt���b$mɴ�ե����Q�0�T��M$���AՀe�W#�v3�k]\��S_�ܥ���p�Kn2�Ut�.`�Z����m8��Gm�3g]��.~��^4ϋ���d2�Os/��X�C�ȓ
��f���\��'qc&�1lC4������6ЈW
M��o�\�9�i��@�o�%K�`ⷵ�HN�"�'ز�{!Ё�Lڍ;}p �/��i�Ah8��x٪�%�߱�D��Р���������hb�7��L?��!5�P]�2��g�%?��������I����� ���4^�.0(����d�%�Y�^@�I��B�����(���w�����Ơ����;&��	2i�%M���޼wCڻ��z��3z����;O��*�@[�]�dL��w)+�U��N����)���Z��|�][)��"}+�>x7�b�h<�`>�3B��I�iv�(&*K!�\?m�)էR�N��ۈ�)	�y��{o�����0�MW�����i�'``?IׯY��D��[G�s)U��.�?-�#����#Q�=�bϨO���t��Y_�R��i��%`����_��4xf쇬��e��=��B<��m�:��KF$���5|�T���^Aɺ4��k?n���ݴhZT7pa(���Oz��3$lś�����
T��
��<��vD�0+4�<��O��FH��o��)�8H9�Ҕ�fbi�M.�Ů�)�t�G�g���+���iJL���	�QzY?����-R	��>kF���"+���@$(��U��n
 �$4��V�������q��Q'x>L��ϚI�;ᴽ�&���f���+v?.t�ɟk_L��(Mhz`/��S��3��Cf��\��N�Y�e�?���1�7�<��^�P�1�b ([(�hF���(�N��S|j9����b���]~9=-��6ÎmV`�`@z�O�_*���_s����vqix�$8$�E�ÿZE�L<�
��a���c�`�b�ȗ�<�abEy��I�%[�hj����LT>{�������8���:P�6����np⎛d���N�po�]A(}�5#`%kg��9P�RIu�F���L�.8�]�E��o�l�R�^����܇9���K���67ͼa�R�(<��3f��pVPF�X�%���>/P䴸?����1��G��� 6��I,JV �)mR�`����S��u�\?�}b�$�9��B��܆�J�燊��)�o���¬�^���sŬ�'9�ιUj��z�x���E��r��#�3q�=t��l��DG�Ma��}�7�}2s2��)e��Qf�O��E��Џ����B��k��E����3=�SWF��Z1�����2�fa%�7-Rg��h�o�GK��� �&��8g���d%�s`yf��F?t�$݅ŹA�m�2�!�|���D�Y�8V�t�w����Qo�>��a�UE͠ŀ$[���n��Y_ �iS%�2_���5Ú�A������*qK�lWf���tpGb������T�%Z�ϣW�/�R�(@ȫ��gIE�jf���	�'���4o�)����[
u�r�6��y�ƾj���41%��=|V[�M���Tv۾�*�o��~�*="�}��
��3�M�/�ω��Cs�Qr.�8G\�W�5�\4� {
�d(�ʒϣ&�+)����+ܭ�N����e�k娽^��UY�3.r��tA��F�
��6vR:��$܂@,� �k���˂��*��K�����@zX�����[�Ci�`�O+���.��@�+ֵ�
�ƙ�p���ނ!���)p�P�/�E{�i?KWx��^y�Ck�	�A�#�Q���K�(�4�+m�Z�1�MF� �'��+�ӹF�ʮ�,(��tgyv�v��>2i���8�-qu��!MlGybY�b�I�յ��:��J�Rv1g�����aG?�J6g�pUv3T}��u���4��H�]����Qmj?0f�! r��>4�G�1>�y��rU�B4�s��r�� `�<������J�kQJUP�.���9���1b�V
�~,� �+tݛ]�]���'�#��E��,�\nה��m���PK&�����3�ƙ�kËx� ;-'�Y�~�ֶ7�[q�	't� 0?���j�߂�Ƚ���#ܔ���,R�����őLI�Ϸ��S�ea,��A���Ϸ�q�(�E9-	����C�O���^(���y�� k�@ G	UKR(�`�`��*g��W�>{�
wXx��jf��JN�0�9f����>���X� .C��!K��t�<o�g��ЋpR��ojXT���������;�H0,���DCǔ;�%���V���㥀��
`\萚S�����A����V�99���`�b`i��E�	��H(;�O�1m�&�X�ؙ���M�+���y����%��V8��<*yI�����wg��l�n�{d7��cǉS�UB����*��?]%��f�Y�׭8jz$f����>��l�K�'�����cOsn8��F�IG��˼�w�рe���uE��m 	�}B�Z<Qbu�Ct�\�3 � ���Q)%�NZjPd��e�dѾ�v9��{�.&���h^"7�2��?t?|}!�����r�Ԋl��&y�����hĠ�M�s�����BE\���sR��ڃ("R�Qz��oD,��ے�E���+�׽�
j�w��-�$G[����5�O!�5������2��?�ON�Ac�ސo��!����i��fE+��!�5O<#%��2o?�_�1K����L���1���P�� Z|��Z�]B�
��	ό��v$����t(e�$��Q��I F��n��t>1����{cd:]����Ú�U8����>�s�6�:���O��iQ��㓳�f+���L��ήzz$��y?/j���J�	�fޱ�n��3�`�f�'DTP�xw�֗3�Ξy$c���%E�~�Y`G���o������{�]�������K;#�v�����T 4k��G�S��=�ǈU�����1�}O}L�(W��a�B�F���o-Ƿ������?A1fKV�ҭ�ΩP��#R��_��֋�T�ʣ�0�aZ��
�(m.�]ϙ�Ck���%劔���yw�5 ���dԽfZF���.�j)� E�j�g�����m8�O�"��fW�b͐�`mP(H��d�{W������3�8����R_\
�əY:�[�j���$�:��W�l�?���o�}]�cW�0�}�7�W��Ώ�%m Ћ�c���LvTy��u��d�)g�=xL��5`E
������j��P�{��!��Q#��!`A�B�W<q���G)Yԉ^L���)jqte�gxm4���@P�����Ƚ`{֣�i�����p�M�$w���h*��Tv�C�>I� X� *#�MiU�� �)3�Sf$`sTr�a�	y���e��fa��K%9�.����nB�뗛�f^��X��A�|͐��ron�2\@4��c0����֜:bY��h��ۅ7� =Ziv�z�����r���{�u��~�����C���
�~��N��u��4c.[��V�u��ʈs��PQ��La��x_g��TG���"a�w�t�w.6������)Q�е���|�8\C%Ӿ��t�/�{��Ns���iB_�W��Ѽ��#߄�\��Dl��z�>~p^6
dX��H��)��E��z����"i#$���z�3R�{�y-K�����O��o_rv���r��ݺ%�������]Z��L}����A�Ovs��ֺg�&��pG��T�#䗁ⰄfE}�x�Oܘj���`��nU�w�0�3�[�ο�*�n�z|�Bn���(�͙mF�J]&	z0=L�2[�MYn��� P˪LV��76�Ѩ�d*2*�>��a�
����3���ȭ�*�@h��6$��L���7���)�"���\7�]u��܇�D����%p��a՘����?۴��Tz�c;/���5���G͖����{~���$5cG8/iEH/����U����'_~K[�kL6�m�q�oĚ~�G�-�R�,��K8Z.�Kmn�0�%�'Z`�P>��dŤ�'���T)��W�p�Z_�H�ꚲ����e��*���w��٩��],֭��ߺ~A�ƺ��,�1�"zX�����c�Ԕ}���Oi��z���C߱�p��`�&o�!�@+fju��U���'!��CϼJ�.������x++�)6���W�Z�W����p@<I�>�/w���A�U���$��D�K <iA���_�i��ӵ &�Rw)�;>�{=P����V�/�@d��E��8V2�,$��%���$S���<nXV��0;��K��J4/,�SL ��/�[�ǟ��2��e����@8�B-$lC�.FE������3�9*���N�%ͭ/ir�!�}�VY2��)���a亿^&R���y�Lw�ΨA�r,�z02�>U͆�u��U@I3��ʢِMB�Wk[GQo����ؕ��	q�OQ<,	y ��G��*�_��^��zgZc��6z9C	<�<�7G��o��yv,(S��!^\4���C�nk\��l40s��XFq��X��[�'ϣ�Bj�i��"3S�	s6���SVˀ��Y3RF��y����X_�;|�������H�}�j E��L0��eP6j	�I�T+�n�xG�9�Ne9��	�9,��<�9�n���h�C��m3�2�芍�x�ĭ��O�B�V�	#�"t�A�+��Z��ki�x[���B���i�pF�����V߄t�(a���x=i�RO���ޞ��<rK#;W�66/L�;��m�ߟ�a%��b�_�ʼ�f��}�!g%x
K)�-�mBI��䭀�K=F^�`,,�������C"��{�6��dH��UP� �|�T���\��0B���o�Ӥ�7썑x���lm�k
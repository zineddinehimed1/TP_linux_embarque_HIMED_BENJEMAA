��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���|���t�9?T�]'�=Ө��B.8��k�����F^yW#��������3�����W�\��U�mI5�#��A��K���A��]�A����?����:*�+!8j����rb�Mm�6��퟇�1��忥VD�,�*��sgI�%�1?���p�hP���8+DE+4��
*��i���� P[:_s��&O���b�������Fu8iZ��>��U3��G��'�2���nq��K�0��P�ou��UDneNNĒ`�'?2�6���Z��}jEt^jH�c�Po��E�NA?��X�̇9}Vf�]������1FRo�[�ch ��*��_�ҳ8� 0��퇛��Ò��PucLԽ����ԙ؂�{햋i��������5�2H$�,���JTѶ@�Zǲ�f���%��0�ޖ�'��F_�A��uf]Y Pq���3<wO���#x'������*�͎Eoa"�G����K�-�Ϲ��4����H�T:��	-N�Hn�M��GY���I�����T� ���A��+�e1�]E񹼷���M��Y��AU'v�b�l�kb�6�a�!G/AJR�xo1Ur;��N��p����&j�ibp�U�&)gP��[��9���zJY�-3}!��MT�Ev�δo(��e&���E�a���uC�E+�v�c1���g���"�YV�
�]|�.�c河Y��ݤ��Y���c23�����r��(��( ��-*���-������n�5]OC����3L0�G�]}�$�̥Uhb���oG.�:��vWAa�F:��S=�R��aە2<���	��N�^W�^H��t,����y�����2%ir�-)���#ʂ�$�k7;��ֿ�'���۬�v���_�ne���[Tm��jD	���?_l��7��T%���2��=ȝWrS��qY�u{�������?�7"�Ipo�H�����8,K��;�r]"��a����{Wk=H�-�R�+��nVJ�� ׅ�GE�@���TW�ѽgg�E�EދC(�����vx:/��r3��Χ�j��H5~_X� ��f��$��ܙ��gI7����4�:���w//�.�I�:��N����s�π:r�m���5�-䳣I��)Jי�>������H �T8лc�%RƢ��	��q�8������P1xpꕆoؗ6��ST��_s(�v������� ��L{� �sA=_���8�U�<$�*��&u/^!ܔ���yHy�6q�x�ʑ�����&"�5���Q�e���4��x�z�;T��8���3�)R�}lae�tY�y���fq<��.*��4>�V���7UC������4;�a�ImN�'�Y:��6+���
��٤_�0E? ܡ��{!𰘵����o��5(��k"��\8Ύ��N1�V@�i�5g��ž-�9+Nח�$��xUj$M	;��P�y�t$��g���aD�-�X�5A���e�l�V\C�{��-��>m㘲�~�{��h���`������0���D�i۲TN����������?Q$+�@��u�	�p�j�l��#��\[	��#�D,�a��.Z��a�O��Lw_ ���!�zjI݉*�r�*U �@eI�Ə3��ǈ/f)�d{aiPu������Sg�4h��=�?W�����9>��s�G��:��V-�^53F21�/ZS�k\W!o�*���l>nK �1L��:����A"w���;�@��O{��>����މ�PNFh�r�g[���DEp��sN����vq,е��r��??�q�Fz��UMR^"�L8�[�3j-��S�6�����ot�ԓ�Kp���_��㷧��W)�Zϥ��7��8�mU�q&�f�8ћ�[.���������~5�?�L��t#o������N�V��Qv���:>4��Q���vGaH#9eAA=�f]��6��8̊NW����W�b]�u�^T^8����e���O�>8�.P߄�mJ�`4�`J�b�����]	�Bb��}��(�L�C�գ"˷��s�NL]���9�n��m,y?V7EO��2��m���T;p@P�����v!kC�y,8�H�}�~O��N�����}�ឩ��x�����f�{h��n����2�6���I˘fX�m�˳F�sd�%o�e��q���J� �_�(�~�����Ko:�^�=�>��!ۍ��B��F?$��(�<��0!)eC�7p���f�e�� Q��s\��S��� � y"y�Xj��e* �֬.�j��AǠD�5�Ʊ��0�C)�	��#D"�G�d��\9O'�d��.�1��X�*�;���sǝi8�I��gS��ؼ��}��Ie!\*�5��Zp'��@�;�n�&$ZN��j�"��萯�ۂxx"�-��I%�Lɏ!�D���b/�b8��5^3{�K3�2���|���6�©���%��Jޅ3�� ��x�[Y2q�n$U��(w���5᥊�¥�=CE��i>7�紪t�NHIiyڃh�n�
�J1��u��I��;*H(�7�d�B�fJL^�fC���Q��q���]����ؙ��]����¹�Ւƀ�.����+k�^��Ä�]x��u�zT'ٱ�d2}9�O���w�S��tWn&�1�o��`�ガ���	v��f=S��c@��R_U�2�0f�U޶%�
�?諂�� ÜO�7�:^�H3�k@a9/:8�Xw�R;��c�۝��Z�:�C�@��p��|S�=�����^�q�7�8}����ه�T��}�|-�+8׈��]��Q.��j�'V=����I���q��������<�d��r��ᇮ"�8�S�����3�Z�^v*P:�s���˔]VH_�tC�\&���c��(��BOK��������8�m���\hp��^��K���:��(9�Es���H�Q&��!��F"�<�]L��t�V�Ȑ�I�ĨF��|�i�����m]:Gb㙿C�����f����R�x@��ö�sM�����k���_�
q5M^b!�7-q/���'�/��@��y�[�����7K�E���G�W/d6��X.����q���B)��Rjot�q.�v���D�q�C���Yٕ%�~��P�@���}�ѫ� �=nu�Z��v��@gL�vFƏKs����eG�\�����[V�S��y�A"��q"���jJ����R�H
�"����t�7d�w��`�p��뎍x�Z5�
�	�)��I�d���1�d"�t�A��*MDԹ_sw?��.ʧ��D�*tq�I2���'�@l���\�b\���w�� �P]��Y��
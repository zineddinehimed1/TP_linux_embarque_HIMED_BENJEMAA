��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���r c�Y�mI�1M�Adb�t,�i���ʂps"����1�BEp�e��mN�Iq)iv�������K�)�W�кn��YcRt�W���$�(��{���h�J��=�:c�W�K
�X=�ېI)�K��F�ź<��ߑm:ti�I�x����Sx���45�8�c���UE�>�yN{-��ޫT�%��#�Z��h������^t�g��YKa���o5dw�ޒ��MD{�����,���<���K�~�5�cS^\P�zW`q���(\������K���� ��E���?�*������+��QY��ܤ��C4�w�E��<Ru��)�o�$,&���8�%͆V��m �]:�%�I���J��Rjy���З�%���b��ԉ��T�d�ו]�Ar���ΩU�-�h�`��c�]��+�V�?��� �&6͜c�^|���SW�2��h��c��%�Ⅼ�\�:r��x���K�1��w.ؾ��$e�-��Q,z�O�d�:75L��a�"��v�4-4@�sl�no�� m�=(r6ZB�*�q��їˡ�h�ZT}[LրYd5��O�<���f�0��ָ�ܪx}�V��8�V�wl<۬�"W.2����->;k���Cx����%f�.v��y>�������/�l���� �[7����?�s6�	��QM����Źi.Ԝ�9�׼P��0ܦ�Q��]S?�%���1醹�q�Y(&><5��"�E��i���ڴ�{/kwK�o����뮄����n��|���}���w��V��(�LGv��M���LBQ�ƶS�]�es���Ƿ���P%�J�c����8�bHgR���	Bej�ƶ ������W^9�uL�B	�$b���烊�PV�wv����j�|���qBň����s��Fyfv��uh�r݆��<}Ǜ}R�;�� ��k��G�tWG��}�7��2�;J�L�5�^KWb�S*��� $���`\�X�Z��`jM������N�ʆmڻ�Nr���T�#�a)|c���1�mDP~ D���W_�6c��b�K�l��!��CjRb5';��E�f��h�1eP�6T��'����yXz��.�U��ap����/����B=����Xh~喽=WB�J�.7���%?��-Ƽ��nw7��.�E�jy8���Vp���\�o��`G��/�l3��XUo~;Q'���T�)U�ɊoB��_������8��譹x�Y��
���
����GB��
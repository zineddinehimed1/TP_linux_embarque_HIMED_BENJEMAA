��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����P�^�Mqap)%t�?�&�Z�K�*���~O��in�ÇZ2���RG����R����k:�H����`�E�m��C�H��Ё�]]ѱO�UFH�Ꚑ�L
��"�0dF	�b5 �A��Q��+�	-�eD�4W!o�� �@G:�� ����Ͽ���˱z9-�n#��V�G~i�u^�L�������;�q�A�~��4�X�-�]Yl?/�Pa�����4ǱT|���G4'O;&�;�o�u���i~t��n���4-BǇ�aM�ݍa�ڗ_�bF�5�����
�s�c�<���w����\�_UN�΀'�D���+�qS�e-����@�\�By@÷�:K���F��W��MV�p'^���w}�#��
�VﱫIT����tL'c�>�F���b`(6$T�j�{���x>!���4f�R�;�'~>P�V���^�-x�v�:F�4�>I���Qn�0-68�jfb,:$�9>�X�y��?��vLr}p$?�Vw Q`h1���M;�qD� 8��_Cá�;!H���ޑ3p>g��;+F���گ$����`�͈��9D�Շ\����RrԎ j�JXږ?zу[@��;	��X�"���F���b:D��4��"�.�*�8��F����"K��rG�Q{�-M�ǡd�O�1	�9�^��қ˛�:d��>��1<�MaP���� ��a�0�j�\ ]�?r�v��œ�S|��A��ݔ`r��ʅ�R8I������-��@�(%!u셺Ħ1�3� ݿ)����>a_@M�2&o�Τoᇌ�3o��c����;�Q�U���{$:*zt�=����J�����ȇ!�S3-'��y���vC���3�!h�Q��O­�5\$6�14�9�2pҜ��v:nN�� k&�E��D.&��t>�
8��hJLz��R�ȅ�:Ѐ������j�D6B�s����i��4���Ţ|�I��6�ZPWy���h���ܪ`衑6;�Ɍ�G����-�=$�(��[�~^h��L��-��=����p�[�Nq�-��~ۢ"�\{u�י'�Ej#�2��p��&��z<�C��eFp�'xz�%؂�p�V�e�5MI��0Œ�?��Fk>n��y�ȹ3]����$��j(oAV��%�c� %�<r�
u��dOk�vʹ��Qh�d�s�@�i?���AB��O#b�Z4 �Tpo��&��p
�&Sbf>���xSIȿJ����g�1�3��-�@���r�r㪫�хG��--�� �ħ��<w�=�� y,����l�����X�/�Ñ�| `^s5��q�ȱ.���U��{��������0���Z�k	���׃1�y+A�i����7,��M��6�|9%3��+�';��)�E�@]�M<k�Ġ:�l�SK�k?���b�w1�"�EܥՃL�P9�B|�
PߏKx-������i[�9�2U���ꉤ�8��&Yq���
��W��`���D:e�|`����ždjH�Yt�Z��A��jT� ��
Q�u���*��sT�|��6�D��Rhv"L�4�=_����6~p��T�Q�B��B� �l�G�������&�l[PŅ2��͚W�p�>��~#p�N/��E��
�t�	TѺB�|PN�֑m��,��4Z�b�E s`�!^�h���n�h�f��(��F����[�1)�ά�єc8K� ���}��50�+��@���>^�Y�Ċ�[c��z/�$�C��#(�y8|��B�Uȁ�%��<csT�a�?���eZj���pJέ���h�C�~�I��q�]9)V=���;d.�evk�%�[CA�C��3�<������Btֲ;�
8�������W�� ݂ %\K�׿�>�qH{��gQ? ���� T�����((l|]s����ٍ�����|˄߽�V����O�2�x�4�LՅ�$��_��a�@��X4��2['��'��!�7�FS?d�ԫ;�1h�~]Bvg��V%�囄��1�cMZ!��|/��滵P�I��rO6�Np2�^��3 ����y2=�
�.np��U��ȼ岇,�����״��E _��~��[��)��I��u[.
�y�2 �ȏ#F��T��cr���}?��JO���I�����G#�<�,�=	졧f�'�� ��-��$/بN��̴��3(�"7Y
ʧ�t�4;N����A�-h���z_�d�
��@m�}�`����p K(�
�g��m>�oN5:�v�Q�X�V��X�[$�Y*��=�2����=sʽD�n���O����3� �@C��x��"�N5}��m�H�%�B��۝���µY�9A�S9��A��w3_�ɌQR�ʊx�_���%��
V[�ǀ��j���0m����%�%��
�fB��߾�g��A���Zd�1.R�����Posm���ڜT�C�����gpY�M^T�c��>S,�/��-pe��?."�pk~���������7z��ǜسw��5�O]Q���N�0��u�"���k�A�_^���0t�\	�y��+��/��
KmQ�Dͳ�h��^ױr��ܢՋ�re]�,�k�����osi�{�j���d�3�<+.L9�����!��7��mɣ{�⛢匉�EŸ�YD�t��_\���F�\�S"��m	�v	�ۮ�F�'��+��^-�;{�����'I��g�s(�^�dLŒ�������$�	oI�Unsm�Q��%�P�쉴ߚ���-��z���@�ێ�{K�X�6J��q���l8���W��Y;�r3O�SSW/V�]�mAhm���y%�P[�c���A��h�0TQ%���X���,�|>:*ա>�(�D�Y�>p��"I�S�����{/�)qa�H_��>�#&���5|blP�
���
���⻽`2����^���4M�aTK:aձ��y�a.���qKU9�ߩ���!����\5nr��p9�}Q����0��Y���5�Y��1s��к�>F�;[�L��+�A���򄩸Z.)��~u<!=����砨2�jM��P�K�?@hg�U�tJ�;��T�*_�Ң�qʮ��;n�^ya��'��GMf��q�����L��+���%ZK���'7�F��'5�t��G<*�XPψd(h���l�b���u����q��l�;��:4�e�T�(�#�^˙���ۢ�_�	��Ի#��D�{ ��&*�1��9�ɀ���"�3p���r<�,Ip��:2=	Z��WȊ�bOE���~�#6��21�.�y�/	��哣 �% *�m5i�S�WO�y�.n���?q�T��VbH�\J9��h�s��yTQ[�l�����=#i�<�,��>�{f:��9��A�Nq�@�%hU��/YSrE�qvoQ��n��|P5���+,�>W9����!�JX@m���!E�[Ko�9o^"�D1'������paN�>��ڑ�� <�zϫIp�Z��}'�PM8����E_g����M�ҽ����5��&��Z�{3�Y���}����QH&S8z�z�|Yg�q��遼�f8%W��-������K�����̫j�n���9oP^���7��޼�sI�ʝ��x�#ީ�VW�U`�W��nWq��ura�đ��/l3�T*�sN�T����	���D�9L�zm�w�Fҕ��~Xe�?�ׯ�mo%u�RxO�Fܴ�G��n�����r
<�X�Ā�s)4�C�&1:n�-}��}�bu�e=;�.�"��54�K�����6�74��gj������W���Ef�J�-���}��$���+��%�t�ѻ�3���B��O�i�QK\�K�.T�4u)��L+S��R���<������<ndp��k�	W���g{JJ�����C�=ՙ
֘��~��΋�L��w1<�>7�9+��jx0��2)�)���|��V�y�r"��I��WYm#�#Q���)�N|�qjB�c
9���$P9\���㯁�*����+���������6�ԫ
�+/��"�+��?��N<�d'�D�H�v���Yj�d
��5ك�`�7�G2�����;	q}p~�/��-A�0����G�l��@ P��`���P�c_B�S��e/=�D؂u&����|�.��Ͱ7��e,I�k�(
`'��9�!R���X�ws~����q�h��:��@������ÓWo�*L�ss���G��$v�@��V$ソǣ��3^�L��9��4��|����|T�"R$���Q^�k+�{���A��8N-!z� 5�)�Z�I0���TK������L%�=�W~\SE����h(mX �7�?n^��6ԛ��n,�4�zULk�S:�	}�'�����1�G�M�m:����l8�P����|FjƢi�n�<"��G���!�IQ�jp�q���4�
F��M(�5�:��E�z�hf�*��E�"8�U�(E׃f� g���,���x��-�"���{z���!���^�-7�����-�^�� ��nO�LO�`wQ�$��qc�P�\��;��o6̬ d���3w:�9���cܘTt`���g���&@��9��Jm���'�b���:K�W�i�<
���m���:����޲ -z)���:j�� �9>�hyY��՝��t���ja��H����f͋h�X�mH5��2-� W�|03����cQ嵝nӃ*ϟDb����:l�h5����N�m�$��#F����C�O�
���4�{�F�'��\�f��/E��Q��yW����aܹyz�/��9�F��sm��ȵ�����N�@	gõ��B.y��-ث�`<�_#ߓ��u�����6�{������P��p���{9�o?����)��7oG����!^��N��=n�Z
����'���b�,]���WK�V�@�$F�ZaIYB[�M,�J��]D�R��~�=D�[���d��*d�lEFA��7h��!�&q-R�0,�j%|�?6��cN�<r�����z�h��/��-�i�yo}��!������Kroi���� ,� �hu5�����O$:�Կ�A'q�U�G4�wt����pjH���U��P.r���1|�ej.6���V�%��>c0� gw��쬘��l\�l�M
��#.��xVc��{x�+�x�S�ѭ����
�a��G|Y��q,/��{kmD"���c�0U���Z�Xp�GR^�l�8'DN!r@��돔��t> ;��a��A�D�����{ʈL�����$?�CJ�/xO_�s��z���f��wˎ+����]�V�=���_���و�w%�DSy��������zC!uK���N���u�a�2���)��W�r�|u���!�M
l��_�&X�hO�:RTt>("��z�:���Y���L��v,�5Q:�Ǧ)ݛ����nf��yJ�;RX��r������q�o����+����M�,(4�;ŋ<8����( vq�V��Z~�C�i�Bą��շ\�Xw�N��m�����E�鐛<&� \G{��f�D��
*]n'<
@�k�,s����d)�f�h�	%-gziҳ`?�)�r���Q�e��
!��r����?�RUX���a�������d��>E�o'D��ex.��B�c�Yiw��}����IYd��F(�Ma���y�e �����������]���}��/�u���-!	-5õ Q�.$�0���̳����(L�tU� �����Aq18qd+�]�t� ,:wZ��2������"���,i�6�L�m5�D���'��~%�j��Np�V���6��m��w���ru��j��}GX�<0�DP��)���dՁ������F�J$+'�pM��������[{��2�c�����3�W���W�Az����I� ۘv���b.Z�R�2�qOɋ���X���NY�zk���i5��Ҹ��-lό+C����_�JʗUy�/�9
���9���ې��jcst#<�N1|L&��]ֳ��gdy��sV����>�C��02����O�r�R�[q=N����~;9�2)~�_��P���e��<8�n���2������/�[{W�&_��j�~�AX;�m�����8il^x7g��"�m㺭�fjpR̂�FW.�*��"�;�2�#��wogS�]y�Q�����k0����$���`�k�lr�h��p������j s&��7��p����@;�u7�V8g��1���N�?����i��_� O��T~%g0�g!Ga�Sub���������	�vP��b/;	m��e���nx�Z��"�U��o��t%A��dw�����:���R��@�����]Pq�E�q��8�]'�S-Qo������KYp��f��6�b�픿Q����g�o��ۚ������;�� ߦ�5�(�4��Z��$A\���?�s�:������sN+6���ɬ���;����;���{�+����/נu�h��v��R| �/���^g�T��(QG�n?A�??�f��'ļ�d~�T�����9�Ң�����]�C�[_�4;�mա��Fi@�=3����M�:��7z��� #g�O����.ty�̛2��Z%78�|��B6�oK�ݓ/$����̀.�Y�0X�"�ԘɈ��"]B�7$z얡����z������d��.~��3M���F<J|Y84!�1���'��Y�$udq�q(�z�TZE�\�.*+��S�W'F�1�;��e�d:��a�o	���I	�f'%>�����8�<<���xdW��W�Z�ٻ��ޖ;{ުR��8�ޛ7`�Ea'8�v)�c>-枻� |T���]�<�L� 9����O=���nV��d5�mBHY)��})Mj�g��4��zE;=Ks*B�8K[���^��g��ʟ�x��(a�PV5�e��1qL{�:Y�P��s�����0?��7���Ã�Z�F<��lJ��+��{�%���\��C�l@&5%�v�ThOI��K�)���Q���=��2�����"��=�{���tקx&��%�B3~��A�l�22�8>�E3`��d�VYz����<���=�ʫ�Fs�%G�};�x�J�jl�Uo��D���$�8��p݅O�ۏ�m�17b��7��p���t����2LM���C��^ߡ��FJXx�/Ds��	��רf�#��2��NB?�،�*n���sD	4��{M���8['�2W��.m�;���[����r��"]3tjo�O$�������|k�����e�+/�*:y�3f����"�����7.
�[%������Q��J�����2��
��ͪ���'j���1��!��L;
�c%�E$Z���#�&;�fL��?�81��;�\�w�'xE�uӈ�0Zw��IvJ��آi�DW��-���ސw�)흊xΊ<��h�N��`�v��_>��n[��@����#���}�[+��y���%�y��dno6��ߟMm��Ū�ή�2\9�m;ݮ�Jo�Cu?VZ[f��H�3�>�otH�K�M.G�Fk1Q��C����1���x�M���*�����B�"b!wDB��6�� �����wEr��WQ���4��!�Z^������5`U�@)*���(�Ȗ�%ʴX�6�I�33��_�hY|��u�I�XӫY�H�}���NZ��Tc#_�AF���#���Vݒ3��;�˦UV�	u<U�Ӟ���5*���3�\�����������B�3�/^���t��5#� 9Gq�j���E�`�ZG?V�zk���Aw]��@��D�e�����@M���ּ���hTh �=\Y4s��9��]�a)i�0�+�i�FQ��b�:P�A��l:�~���H��:%/�s�9���ǐ�j�Z��]To��z��w0I��V7�kK�N �-�|�{h�&/Vؒ�~��r�	R�6�~~m|6��ȍt�A�>RZ~x|�5�&O\8O-n�>'�垀Y�3��I�$̜Q��ң��bCkh�2)�Wl:�*�p<!OmR�
�^�NDB��z-�qK'j�]�����(�v��Q^�s�Ț�� 	��a+�t~m�
���Z��q�+R�ilyl6H4�~��N�NO`��q6�j��D:�5m�L�P)1m�P�F<��VE)�f���i#��y�����/W_ �L��둒��6-�{o��	/U�zv���f٘�uU��J���a-��qm�屎�2ē�J7��r�5�^���&^�\6��|��o�Ɇ�8V��x���5��V�}����Љ�����ӡw���ߝgTP��C�6f̨���zS~(�.��[W>c�����h����?SA��h�϶����iW۴�i��P�k�/�p6���=���ͅ��N��]�XM&dW;�|p|���E��REP�����:іO��z�YS{འ��3�Q#%ob{0�����c6%�_!�6��<��
V!���銉z���c�����i�E8���4�ec�:MS����7�xUal���=�AvJ���_������B�e"gVu�0ow�S���p S�,�S�!K�A޹`��6���92S�%{̶�������w_s�،J�4�����k����2b ��&k�f]N��{��at۽�$�'X�y���y�g��>C��'0W��>q����qr�r��C�꺭���eUE�^���yt�|F��H��,wn�;��	����H��c*����T������!aA9㵑���;���iQ�A�V0�!V�/&��a�$�Z�I~9j�&�=E�E[un�7�:��v
tY�nl̊nO�.��K�o����S�`���-�*-�����UI �����n>��έ�'�#��*&/�O*B��h)B;���W���'�pƜ`��*��I��Pue�����K���tP5�i�_��Ų.�c��=s��Z��U=�P���7ţ�.���^�2�5����q����R9�N�����E;ƣ���0�N���m�X� ��ۼW[��{�PD�z�(g�dU�t�9��!c,�.��ח��ѕ������O�,{ۆ�w��KA�����s׌1�����<؁;�@�����T�0g�f4�S����s$��<�!Xnb�\�[���\h��ϊĩq��3�݃��=�֚���2�+}�	c����u�m�a@�o�,����3ݞ�̥�c�C��X�+���4[w;x۴3�c����Z�&ϟ=b� _=&��¥Y/��Ew��6��8 �fK�m�Sͧ���]~N��(�@
�'/8^��L��L�Su��#c9��e�ky��	d����V5�`�h�W������ݷ9+b�"|�}���+t�0�@ǅ��X[(:z���c`���̂��Cu�z���)�&Nl-�C�d����F��(l��{�%4���VU��DkRD�A�΄T/���4���|��b6y�V���8m�����`��j.�Y��3�H��n9$�b�PC_�d��5����uH�ꩋH!��p���B���i�hf������4��#5���Sr�h-~�C���{W� Z�N���!���bn���ř>�N�O��i�tثB�ģ����#�l�N� X�}�J�`��t0N�2�ի<�dVq�<W�>��P�m��\EA��?���R�V����u_��*IB&�,j����γ� B�95�i���23!C�]e�����dl��6��!!p��6���m4�����^,��@��o+��#�I���A��ư��
�x���&���h�a0�M=e����v��t3l�%l�'u�(��>�BxW�
޴cc�H��z<p��q��T��:��6GD�;�m�f��"���p���!~�8O��%hTՑ��@��w�E�<�Գ{��%��8�������1�^>/<���%O,Ӯ��/��I�M(kh;�;�ջ�na�� s��g�ۡL��n�.�{�$���D���F׳��~0��$�<��?h�O���[{Ye;���r��}�O	�4�F�pW("l&���!#y��>�<#kd�{��e[���V?H�~I-X�!���W�Y ��$�'�<\�F��� �S
�T'K:p������z��P�[�:���]�.g�_��%21���메6Ж[E��{�z�L�W���I�\I�M-=#�7z��}�K�bA��O�����S�S�6ce���:�rߓ�z� <��e�R�W��m鲌�<�a�d�>c�U���šq�k����vÈO�x&1��H�̺�0+�4P
'���c!j�E߉=�y�GP�k��s2��_(aNO_M���0�#�g�9���Pf�Q�iK�A�c&c�^'� �3p���QX_z�����B�o;R�V�9�l��ga���N�����&�Է��O��Z������"�gߵv3w\����^h�	���K���9!7%S�neG͵,�(��+�Ud���{LW�(�җB����A}�=��}�@��`<HI�� v�L)Xβg���Ձ�MS,M������%�3& ���O�n}@_xyeAr����9b�dpX���4�9�Qd(��I_w��8�"$��x>�v�1�ޔ��xZ��<%������0I������3ݾ܇��h�����r��˄o�ֺ���{�Ʃ���-����󬡃�WR���E�Tf��3�����T_.�m�$�De/O���I�(!ڏN�BF0�w�@f��@�{�a�E[�aL����G��;-�������3P؉�wɩ!��F�Ϋj�4��sxN��gWÎ��U��cH�%��j_��M�v����P&���U�����t$��E�/�
�xd-Y�p?�8hv�QO�I��0H������&r0i��K\��Ѯ�si�YálN�D��4��Sщ@:���Aļ7;�f`wk�_�-M��?o@*[C6�qTˏ����ˋ��IWل�����MdP���3��}އE6�s��V�����\��(�X�ɟ��)�*� ���M�Ym�h�kp�� �^��叽k��QCLJ�̭�-g )�i�Γ2�&M{(z��G o�c�R
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��׶8۞�@�\ږwiܕÜ��=r(ro�fC�pr�L�O�q����6�|��3�Y�	��9t�1�HKjQi�i�vE��{�+Դ	��J6nsE��739������w����׼y��E�FX3	O�O-b_;/-P^@�s�{x�y�rR�%�9��\�Ÿ��ƙ"K�̄A���f;����29������Q<(%��z��/4�f�Q��`���4Q��g���(����H�I[K��:wO{̰�覣�tfh��v�]hx��r�N������EO��a���2���N��Y�2��6�U���R�X�P�(SI��ӵ�͔�-#�'j�(��uK����s��pиl&2R
�E虩�m��l>�f�J�=֧���N�~����zõ1kѻV9��g�19����b@[�75����)1�c!4�-��`�yqU��:�Dڡ�]#��8Ba�Dd�h2��v�oR�L[�����֭�cf�f�<��9�sۤ��!ٻh�t)�A(�9-d���E� zd�OT1!�j>z�륯#r%�K=��ȹ���K�{�/�,PD%�=ˣ:W4���M12��S����V[h������{����_-q�U�����?�lC����v���1�X�,��SJ�Pp����|�T�����.!�Zv�0����l�>۾u Q.A��k�������	�0ox���R��`��+���;��tEi��h����JIg�A�}braeM��r��K��@���X�S�'��Y�-_GC��HŠ�� ���6* X��o�N���]g�������
3z�� U�e�@.�n�;�E�*����?���PvV��?$� eR�owم��9����78���u�I���b[������&����W'^4��$��s�F�l��O�n��a��d �����<SӰݸ����.7KF��2¶�ݲ\@����t�/�fA�[|�Jd����"E�A�=���AD<�4,K<+̑��>KA1l��ٵ�͙/�}��������(|��1���pV揔QQԉ,�o�k��N����_	|�8�p�<��_��'c��8-'��C<.Wi�^��v�������&��F��M�z�����Af��>�t��4~l�bAZ@�c�@���t����]r^��]0�˄���T(ݯ�`�2 [�?�?3r�Ӽ�����੆���O��8�U�y�%�+��9'���j�j�E9z�/r@�s��lY�+ gĊ��f�^j����!FmYh��"Ri]�n$33Q��o��ĉ�q4Z���9��:(NU\�_��;�alȝ�ߣ���ܪ�)5;!�&ҫ�����h�<�R-}�ŘC�V��U9�֩��O�sZ�H	�1���w\j�S�b:G<O���Hw\��?�~J�0]��x���^q3+x��!��[���=O����ݴ�jDo7�;�x�o�Kua���0�29X8?�qXU.!�@�E?[ߞ�|�f�=�#��Fh��#�U�w�b��ո���⢱�?���`' =���2r��g<�V��:��[<��6\E;va۝
���/!��q 9~�¬�)�(�|`�K��S넰Q#��<���]l���f.�p�U���$׼�
J/�L�>���W��Z��<m�G��a�zɎ��<��ĳ���Κ����)�xB[@��@ƒ�]f�p��.�hX�]��Z�o��������LL�5ֳ�OFܙ��b��H��h�n���ǐR��yQ>��D]��-���d�5i��
F�0���
Ɂ���΍T�X{IfU�	љ��A�"M|��&�`޺:���1qb�]�{KC�"*E5�ΛhS|�������0�`��)���kKɴ��d%~:�Ņ�Z���٥=�/�����8ᔧJǨPQ�$���]�|����j~Jd�4/�⛝�=R�oba-;?�	/C�r,�y��|˯S����E`��h���QL%����Baoh�p�� f{^ڤC[��������^<�	r`򓾊�-��E�;�z�q��ޡk�`����{lz��X-�}~&c-�!�j�[czV<.���0l<�<�m^�k�]�-ߌ���WR��
ݸ+�,���`2?^98t�Vy����5�siת���q�����9�hu5����E�f��An' B�E���E�b5k��6Ф�����삶��]v��2:,���q����͉IW�LǇ�Z-:Hc
?��ы�_
�V$;�w&�'�'G�D��4r=�pT��c��7{it��B��?���R �|�"ʓ/x�jLv\�Z�[X�S��9�uׂ*���_��:;�7 ����yӍ��+O`R�m����~ի\����o�����uss��4e�/G�����7���E�@��e h]�[��f��00�Q�u�1�*��$�"�|�$�����T6qv9�8fk屏�d�ig���qan
���������Ki��;�ϕ䶳���	�����wڀ�|�XF��S���?FkB/��>��CNP���Fo�Q�z�@��Ě�)��q
@��Np������tT[·���U;��zH9���=��ȩ>�����ve�4AJ�C��@���������ߍ�sC;#��V�	3�'�0+� q.	u�<�Ӡ�4��>���/�4�]��_�~�JY����GU��"�Ky��e3�Dn��k.��D�J;��E��vsĂ(�a%�y�?B���%�ϐYt�Bl�o_؁���oUuM��7�8�"���0j]Kn��[�4_u�����+�bJc�2�!DHJ��ChWM��M�6A��N��9�=��,�2_[:p��}1Iܧv�f�z�Q��w*W�y�d���j��ɿB�F{u�IeD�r�	��?���r���(,B(XrM�Δ�2}�w�e���HB'��E}he�3Jߑux�{)�84��P4�D'�<ڄCn�����r\�]L���G�Zg+���4�ęF�T�'��C?w�'}��v�M�.��ɪ�T�#צ|��ʛ���U �� ��9�u ^��1�?QԼ�� E�@�r��j�w+F��d���~�T!�_US���.� ��E��c�A�]	Q7�S�� u�/����=�,O>;1�!��%��W*$s���SS���l��zP魕��5�2�%eO{��pTA�U�T�2=;�S{�hq�h�j�);�M���56{v��:V��|z� ���'���AukI��c��A��Kl��ֱɁ���5���_����s,e��7G���Fۖ� s7�}T�I�s8��U&א��e���^1#��Vb�:8��0d/�p8�ȹgv��������ŏ7���!G�z�"PAyR�Z4����P ��N�����㏑����+/{����}�w��w�s		C`��>��`�G� ]d�_���S�E�6��j�vN�[�MM���9y͙�+�i��\��,xS�U��s'��ԗWf7��IW������8�qmqP��Y`�V(�_7b>wҗ���!<���0���}1\��"}B\̈׶v�BG��푅NrII��� #y0t�cyvҴM � 
�\�1����VQ?�˨�%�ݑ��ہ:#U���Z����F��p�t�Q��pp����W���P����(�p��c��;�$�l^9[^��mb6�K�����w`S�F��ZV�U6�+V�N:~6��/O�,������Mrp�~Ħ5ﵝ���}�� �Z��9�|b�|͸���J��������ɕGYR���纟۔؂ަ1��L����Mqc1v**m!��|d����9�9fم<گJ���g���qg%q��@SJ�!v�Y��n�ʱq} ]�,��V�&�oxش5�Τ��\���p#�c�︒M�gh��q^W�u�����,.�cu��1&}���}��¬ ؾ�[��@��$e�1���#t�<��I.�i�w�ȿ_�5W�L��%lS�GE3��VG����Ȯ2��9����N��_���k�D�oXyKP ���z��<�:s�5��kNƣ�傴fm[9׽StFت�!~��
�$	fM�6J�=����ǣ��+ �=	%y�<��FX?����T���l��
�� �d���	Q�"��no_��Vx�g^��� ���]�w�a�d�j�4�O�p>�K�����h���F>{�L�1 ̨�y�R�Ƴ���\jǧ�1WΨ���<]� ڢ���u����#����-����C޸�]����9SM����#^�m:QF��%ЎvI���x��9큞��0����_n�;����ZǑ|��S�M��ِ��]��ׂ#��Sh���PF�^ e�c`W���������)j9�0j�ϒg��tի6�y`�9���b�_y.6<�ԃ�H6SHi�w崯��k֣�gT!G���0:ν��a\5���3z[�L��Զl�� ��.4k�n�pQ�:"$�?��\��q2�U���q<Qs
3���2\��*K�'�v�����6�`5sF��oN���f4��TX�sEp� ���$&�kY8p�N��Ý
��EdO�Qg����+�ab�F�Ў���@���� �0.�f(Q�\�'J��+N�k�
�e<_��4hg>~ct P�B}dd�.�(6����o[n�E�z#(�a�ӳQe�k�/*�uw9@c) �U�uɏ�Z�y���L'�Pq<��?Fxr�X6���Mf�r��Sx�a�7�ɐ��͊K����0w�J.G��P��W��x�9�#*r������JX�+��@:!Cܳ9�_Z����]<���b���\��k���
�ӴLޫ��[5��De���'�����A��nMQl�r�&\jZ�D��?�N
�^����Җ��7#��lh�����UkϯV}úZ�����Q��a�
\���s�,��a���VJQ��4�8�	D�l�� 7P$j���T����LE�L��c�Jj����Th�����a���$1ކU���Uu}�N,kl 	���Κ� =33���N�.'��eM~^�-t *_!.�MV�!./0�H�}��^�?>RF��}���$��2�?�/�֔l�.�2S�lN�w����h|����������,s�J��,�+C.��X/h8nZ�)������ӥG�����D���S���s��*!2椵#3K׋�q���5���PDs@L|���q�C6����M�m�U�b����#8����-!V��:���D}�o�l[<s��ͰPkJ?�_�E<���QUou�]��ٖ���ؾ�z ?�<׋�p1�x�������(0�����R���g�@�}nϯ��4�,ZB�)����vɿ�4V}�X�г�y���[��@�,%*����
*֓P�`61�/�*���2�C�-w����3|�n��Ꮎ8�B��|������ZD�M����tZ� WI��A�����r�&�";'��#�fK�~#�E$���ݐC�����D�~�LZ |
f����0�~[#OU�F3R~���y�P�+r�
�OKRd;x�����Q:CA���{Ex�^͆�6�O��ָ�l�/� ����b�󙕏M�+��Ҩ��UV��3g�2QKD���6~>.�z�ݺE��8��6箬K& B3͑�mg^�����,d�?h6�0�-��r��~_��ȴ�Q�a���;�-�}T'���*��D��1kv2� }��db�f�h~�UBZ5�6�_>I2KQ�������?���;͒�Z\o&������wۀ�eۮVԡ���T'Y]��J�;�Pyi���z}���r�n��9;:	�?S�&z��yb�å�Dk�Pz�S]���pL�'̚�i��+�����HO��n�N[��
w�K�v�?{m�.�O2<󛱇����P1�f�  8�X.�TpU0�ۘ!С-��r���E�{!�2
H��1����nKya(��E�M~���X��c
NJGF�d�P,c*�/	L�ZL`S"�Ȯ  �"iʦe����Us����k�߻N�ld�g��������p+�m��b��H,������ϡ�i�:��v21�d$�ɕ刜�/u#Lw���x�-����NvJ��اӐ�zߒ�<V��*1�B�8�CԒFD����]W46�@���9;�F��u#خ��y}���t�RcMX���4N��E�О�~���8 ��W<׾�����&^�)�_�p����{����1�ڐ�,{kl�{ӂCGN���<��j@cv}@B���&o��wJ���j�}P
�zZ<����ۆ0�:)���f{l���>q�!��C�1`���ʩ֫�0J��P��Nlw�_byܽ�E
oٔT��bQ��	Ox6��#�љ!�j02����q�ɑ�v� ��̻0�bt�:�gmZ3'�l�y}q�\~	M�r�D��ئ�X?""�KB�+ݘ�p��!O�1[�fWRޓ�$`��+�=}+�X�@�y-Ur�9$ӱ�0-QH�'���O���vG�U_�d�E\˫����ð W��-?���󏿯�7\��:�0�u=��e@�P��UmR*�H}*����f���~��_�q�<K����Q������pU �� ��`���}qc��3�������'tpo<��B_�C�P����?�>��"N)��i���e0�5�dI��]W�m@�M;-�N��~���6ܑf�M���eD4 ��y�^dq�`U�[i%Qt�V,'E� �:s8��$U���?h�bp��R�J:@dJ'LI}n;�nQ%�[}$��y'�H�[
{Vh�*e�t��k���Џ���:,5Q*�)��Z�g葊@|��hÿW`���E�ࡤ��>�C^�(1j����`���0��0�w�ᛸ�W����1YqQM�Ӯ� "8.Lek����Zj��[�u�Nt�R{;�4q����KY �H��,���u��ݗ,,�`@KzQp���d "���{坺ß#>�|�[Uv�aKb�e|N��"���ٽ' ��l[s՘�&O� Q�Z��"I���ef�lg5$�(�񗹮�dfB�2x 
S�盧ш��Pkr�媹�=�w��APi���Wt"�Sp�I-@F��Y:���W�>�>��4��]�m��z��1X_=�	*rs��F��dE�=�x{[�ȡb�yd\^ѱӵ�)���n�52��Ȼ�-��]�p��IMеc�Zζ[K?�����<��� )%�0a���I<�B��.����#������5{�PL98�(��\wC��V,�ͤq��#��$#������1�g�Z�D~�J?E��,� �����K��}���4�r�xʎL����"go-%�2�q�q<�l�6���>ɣS����/��^n%J�W�q��w�:	�:�4*) c�����i�e�䐫H� o����|>���OjT!�)���}��p%�������>�U�~�^]��!x��n#��H��j>r��|-��t,ݳ��!=I�
��K������8ùR�����l?�"K:��IJC��dr�ۡb&%�e��Xޗ�D����*�X�H��p=��$�"?�Jt����n�N���7Y���f�6j�O4��L��ߚOlՁOiW�~�.%.���ꆃ<(ʪ~N28:LX����:ʒ.-�t9��"�t��ʨI�MޤC���H�����)�JT��׭�@4�*��ۡ�]s;��i}��oU.�d�_$ړr�c�H�i��\��!o������c"ɺ�K�{��Y�t�?��텭a��c���H4pO��bZT��Fy=>0O�$���1"j#�oυ�~�<�5���	��͌�$��q6	�����e�bD�!yV*7����X�k3��`��2]�!��e�a fǛq��������O#od�/`�l~�y#	�"/�]��3�Iǽ\;{���D!�zFc���'1�t �����"�(�����Z�?�;z\�%���(K�dV֠�<-D��z�:$�ŬIgVh�@q��V�G�$\�K���gE&��/�^,�T������m�"�R�Ð��	�{��6���F�Д8'"��~pMZ��9�)����s�B��I��(;�{Α1�>�߲��d }1���r�ne'uo3��
�=����[�z��;$"g|�L�I�Q܄»��q�ȹ�,�_�W�L���Ftt2� ��W)�$}ۊ�!�v�o�qC�'k��-��Q�Y��A���9��dt�Z��^��ܮZ�"!Y�?�ԛI;]�S���)>�pc�n	�֚:��u$8����W�a�ɭ6�����ῲ��U	�vh�����$"가�m)J�EtۡC�ԡT�?��,.�m-8?�9B}8���v�P����S��	�8!�{�{V��9h�F�I���2��������~x�c�@�ȱ�}7��W���u��x��]�߹(A�����Dt�`�8���%��~�oFO�UH6pS��������M�o.����Q9B�-��u���o�K� ?ߪ-�4vh]��GP�&�"�&`��0(W�[G ��o��z���ej�����>���2i��cv2R�{�����E�d��$��&�؟�h�ޠ���A[�J`8�X��T�kg��f��� [��kP�Wg��V����Ɵ#����������g_yU�g~Cc�"7����O�о�����u��|u�M߫��S܍�Ր�^3�Zo�L%�F�ôW��p�����n�lk
T8��Jퟑ0�O�����Op�"�''�F[	�Y����j��tc�����1&X����{����0=�^�F����0��������8AMñ�{&��{QЯ�'�j ���wH&��Jk/�P�_�"�1$���EC�`<b-RwkY��'�ԅ�z�$C�]]T��8�!���ہ���h�?�&�?�D+W�6i�U��{t�= V���]�	o��"F�	QpJ��6��ah�O����D�����T3�����8v}j6~��y �}�6</�J^GC��[;z��i:ԙ�����|����[
KY��37����j]�G�C"s^T6��IzO=�d+�!��h�����X�2R��v�[�#ǰN���;U�FT��
B2W=���,,��*�q��O�!��z'����.BX���W�,���4�r�.���7l2m��=����Ɯxk0����ZɃ��UM#R��О��Ÿ~B&g�Y3JN
u'�U:���N_��bFCV���;���R�X(�;V昮�m/	�/�"�_훲M���=��/H$�e<_(����v�i��՘��;���]]KQ{�@3�>6��e�0҈Ϸ�������~��k���v�5�ɐ^�Dx�J��r9�v�>��	��y��᧊P�q�ozz $
���.e��n��fH��rc�Jr6BG��Qz�B��i&�L#=�s�8�6�R��NH�f���OE�O��P��49�aUW[��㛫3eO�_�}�P�=+K*l�;�/(��I겛. ����}(m8��xş�C�6�YB_B����*�9qSX�p9��wX�#�96U��_�q�1�X��2¥H�ME� ���ߌ	���V(W繡�-R�7դ��X�4�1�8u���T��;c��'t(���ǵĦ��[;�b�G��@A�����1���c[�#
�S�	x�,J%U�d[^ ic:�-ENI��6���(�L�BÝ�����([~Yo�Y�$���s5�?��T>)��ʣ#�F�{�����|�֛���u[zi��4ݾ�2�F*�����r���^�ɕ�+i�	5��x�l�C�Ga{�>(�ˁ�8��Q�w��!�����鮓Z)��sG���¯��D��Z���{!�`b�f@�H��Y�H��L<u�#Q�� |�)��[c/|}VDB,�����7�nG�e��F��FR���;"��0J�V�&�>��`w���\I�`ƹ���iҟ�>At� ��Z����N��Ӷx�Ë���8���U�*��8���,�C�9��N%�b��N��O�>UyN���W}#Tu�d*IͰ8zt@���EG�H�њ'�FV��	QQe+�����GkF�
�h���ICT�:��$<_4=*d�������u �4~1�㡊��J���5Ø�V?�:�^K5�3�aUqHW�N��)̯J�߽)4�@:l ���}��H����2�i��ˈ,k�8 ]�tNx�V`�Nő,[b�+��h��k|�Vq�M�Ŵ����0���y�}]����
P���w��V��}3�<��c�V� nX�z{̽���d ��zJGD�5��&g$KZ0G����
_I�����e[>�V��E�g%5C�vT����m�5�_vj� vU\��ư�Q�L�5����hQ�ׅ�Lu� ,~�x<\���a�\�����O3�/��7S� ����n���n��w�C����:�;�8Jg���@�{����H���h����7�u� 椿�Gܾ@����W`k�$��Uz��=L�l�W�q_϶O!��W�-tVB���A6 �6�Pl����(o��ڇT޺z?���W)	z!s�x &�6��QpSw#ra��ڵ��W`2���R�A���)!K�_��{KH� ����R�gX!�v��/ 4s���M,��*�&/	�-���4tH�_�dqX��|U����1L���d����4u{1*����_�����Ã� %~Z����G�����uKC5>6Ѩe����QD Ra��'r �.���	���C�&L7��F��7c���._��ڕ���j+����������D.-A�ˢq�&o{���,k���m��v�_*��`�����sF ��x����m������7���1�b�Զ�t#����P��0��1R.Ns.mꦆ��������M�%H�������(��A�iF���W�27���>��G�0~S\ߴ�O̔���q�>�Y�C�kgA�&����%:��9K-$%ͥPXPi��-��o,x�О_	�K�eiϬ4�Hɴ��q�s�tK��F����,���杄�6���Gk蝽y`���\�6��}�5�^Q�:ma�z�Ź�gНD��MIv�� j�^_t���Ps��T�c[��*���HĈ��O�B  
���]��I��}�{Ɏ)�6��h֥�L�ؑ������Ym�]PȖ�\$#�w��`���P1�א���Z�;�&�Q(0�ta�"��٩�3	��RC��P�|��s�q:=�N�� Pl&Q/Ӣ.�K�Ss�42�1,��r�A�����n�Q�`���ilV&"�EξHsO��~������Ƈ")I������aI2eng���ތ�cYU�/�0�r�@�p��(:�����q>D��F��R~b�|d4� bz��t�@���l��@�PD]�j}�#�}mL3
=X���"�p^�
.#)((���N,���\:}�N��=�xK�,�_jlv��ꧩ�?�/I�8S�����'�TfQ�h�����o	iFOOb�<���������?_i�����P�g���r�2��K��UBm�
�2#A�$���t�w�@)���i�HB萹�,����K
���O�,�g������ڸ�'g-�"�-�d$P�Ե�`pxex��0"��E�OO� ��/�
���S� �C��T=��E	� �}s��H���j�dQ>��zj������L��ɕf���H>��q��^4%Cj>���1�q����,�wk/�U�{���"O��?�f�r�ˁ>F�?�[�ϣ�����>~RjP�G蓜���� �kQ��@ǳ��������e.��@Ȋ{mӧd��%��cm��Cb�
Q2qze��j��(re>o��[;PB��G�b=+�C]��o!�������$���%w�T3��hOe���Rt��ٛ��泚$�����vW1�h�6���/�C�z���v��t���e��4��5�1/�,�M@p?��
��(�ꃈ����k�a~v	W��Bơ�Y���VZJSD��z1�# v�I��ѐ��m���"��g�]J۫�@������'�"����#�����@�G�V��@�"��7A�*ѿ6I��X��TU#��2�
Sk���B�3 ��fv�,�ǽ y��u���E�`�e�0%D�bb�� ���P��3K��mjbB|��o�B"����54���t�S��k'*c�Y���7~�Wd)��W�H��e-��&�++=��J�YD���J����Ɛ����|8�2�p �蒂>`�I�NiЋ�o��V�a3��(�z
�Tw�h���7EPӷ�wO���r��gILa�1�^bKX0m��|<V�����ְ�h���젋������ic8�a�ū�Ӈg�5>��iI�7�-:Q8���ЉTjI�c6�e7�2E1�<
d���
O�Z�_H?i��H����4���BzB���ĥ^\�I-�$����#H��$���|��4�_]![�d"=���u�6ʗ�(��T�-��Ͳ6��p�L��`u?����SWge ��W��a��y {�(@�\�Z�����	9��G�@��Y�`���g��\��:�d���
���:� X�:�����d"k^����%T���u뮤��H�P&~N� �B�#]�f�]�Wr�(���~��DW1?Md g�5��~]�/���;a L���$3�Ǆ��O��?Q���^��R���]��SLFF��4��[���f��Z���(���d@�49���j}nn��E2�� ��O���T$��E|��CD���F?c�u�;B^�?Cmt�R��f��S�Iw�'����p��8�A#RC1c���YI;*=���=�E��Z�a���T	�!,����=�(0ѺYvy���
��;���Dy��N��ǵ��v�E��C\_<@�kv��Y��S�8�K�St�ٿ�sRB���<'h�c8X W�����];~��Qj�ޑ�ۼi=t~�$mg �����] ~G�W��tj�o3�yr�+H����CR�9ýÅ�w<GF�p�v�]�!5���k���O���ie����>�RSQ�mW�"V�P��P�]�aGr��(Gk#��#Gx��(~ ;-�!�iA�O� q�`s�q׷s���檢O �
��[ġ�7V�ܖ���w�����"�r���o��vhu8�z3yFI"�*�{��g��[�Q�_g��׮�>;�{4#�T��|o{�2� �)���9�P�W�7���>�dۿ���l�u0��i��g,bwۣVK;��E���ݖ��sś��d��{�O.f8^;�4K��loed� �(V�8������]��ɍ���b�{�2������]�ؘS�����]���k��a>�C�:luuk!˯X��I�Ct�U��N�_?�	)��+!�z/��J���������o�R���0�V�� ��C)1�$��#�:B��h�j27v%F��C^^{!���j?��7xV��Xq4y��7`
m�l!���WL$��iD�AW�A����0|�����t��'`�Xl�f�fR����a&�E ��/�s�`�.�랑��jȠ���ϲ�>�NQ�n��?D�M����q;\B�ڒi���|��'7siɟYf "o�;+��
PU=Fd���O 7g���2%��G䕀�t�
A�L�%)}����	?�PH���M(�L@W8da�1[�&������a��� �}(���8����=�/ѵ��;ҭ�����ݠ�@e��P�n�.�j�cx��фRyF�:���=�U҅�=�F�X�1`06������Kl���J�o�����޸��*
���20' K�)��5�����Έf���4���+�=#����Z���
��V#�zE��{z�}Ώ�荵��)�L�7!��C�4M�ɇ\p
$b[b>Uu(�o"r� ��[nW�r�w=�>�O�aw�� ���B�x��ڜY�sY����Aa].���*͈��ۄ�@r=���NdF�k}��<�^�{O�;ɳJ�����]1(cq���ٺ�z�Ļs�R����1��<׀�N>~K���)��b5�������nT�?2d_W�؝����'P-ч|�*��g��rJ���$�^T<H@���;�|�º&�>��I���]Ac���0ω�mq��SYP�΄���;h�i�n4��Y���'����{i�0� �F��u{j�0� �Jh��Ȼ��.A�
5	b%b�ث8_���;V<IW���?��Ā_&�˞zj�Ɓ���ևc�i@FW�W_85�N6<�7�����m�"%�tv{bDM�n����%���jbK4��R髟{����s�Q!R&�.�������ɹu/�k�P���{�p_��.��@>�Áݻ�˃L��~��P��^%zJ74�[<��[�^�vn��\������dF��~��B���_>R.��Ѿ��K�ۙ�����0^;l�%:�3d$	 nyZ�#Bc��0=s"�73g�cMB���#DP0�*��&�bQ'�6��^��u5��oA��X�f<�bxԽr�C�����QN"���CD�݉�*]<��7���x#��R8����劥�f����ǭT3��*����3Ƕ�gˁ�n]$ɇ���K�� J����P�bJ��o*?��x�����Q�p�TL^4���x
�|�+tl���G�\[F6��xg���
�.�3oKȻn�^?��М��˓�z}~;z��:�����.��h�$*�0o5,e����.�k%�T�yz�H��W�q�z@onG/�F'�Z�nӱL��,�<�r�Yn�\�ߘƜ�*Lr�5�8�H��u�o%�7u�4�,�0��CW����*���Z�=Jhsb�Z�R�Șe�!Ȯ��{�m�L�,YL��J�H��~֥�d����$��K�G��ފ5��ۤFM,�Hbe*�� ك�ô�	�`�@����P�ŎO%���^�p� ��!���|��-�IO�n�m��W�i	��=��2�Hת���}='���) [�6<����r���{�P�2<��l��KcYo>��-µ*SH��y�o�����WR��\\�ށ��||����b/|���'�G�x�qY+0>7Y)�[��{"�͑��W���̧aJ��}�"�1�s@��*�hoP����џ��ǻT��oǊx2��6$g��Z]�T�ٓo�i��Ӿf�bT�<r��n�E��z�*6�뀗��>���_�0,�KP������-�e�sj~�]q0���&y�ā���[#��VN�O�u�z�A u�Pu�:�� ���Q�ox�}/Tm����a�dc�_k��f�(�r].ծ9X�m�v*㝨��wBU	F[���c������ۄ%�qGZ-�:�jA����׳'�G�ۊ	85F� <9���J�v-��yMn4M���J�Ċ���u8��V<d7�#J�tՂ����h׬ �B��|v8��W��o��9�o��F\��?�<������#��{���݅����V�k}�4����Ci�3��Lj���d�T���/!8!�֐I�ݰ��lt�PRƥ�a���$3�0&�4��ު&�N�OBI1p23	q0��!��yY�
Z�����J�������$:Ao�-�Pc,]o�Bf�%j(�~O��t����yp�t��Tc�Ņ\�4ѧKh��8#r#�9���Xq`I�%���-PtR��"4]�w��H�"�.���Yў[&�>�;���."/D���M�Ù�(aXPZ�&��m�C3+�Qt��,�Ɯ`�B6���G%�R�=��Ȗ�@1#����m�|����aO|�=��u��;B����U�퀤����*>�a����(}C�EŔ}<m����9����ž	BӢo��k��������*v��t:�o p�y4��e$B�xޝ�� al�h���5�ϦA��T�^Jb3M�K@:;�Ӯ
�K%��t[�/�:��	A���� ��[֨��o0���H�B���]5*��%�,XSN%�~�^��O̚���vv��[�n�|�3��J �[��@���H�����S��>�ʟ�ֺ�g ��}�.��Y}��H�O�{ˡ=��Pa��[J{�r�7#-rP*����V���9�k8�9���ᷮ��u�o��)}�S�=S���v����p3���/mڇ/���	jA96�@^�u���[�QV�s���S���!�S)�g��*C�9S]��-�:I�<ߥ��s����ZV�$�R�?�C��`w35�e�i]�F�uk�G��Z:q�`����x�s*:�Ch0���I�n��Ow�@��oP�=�1ӽ�&��o�]M>T>	�� �F�����u����x͇��h1ق^;���|���&���c(4�߯qN�����.;���a����,8LȒ�$�^+_�Y��{q'H�	jҗVe�`꺼��%ߘf�cQ���ȩ"���� Q���-�r�5��	i�+Ł��s��mv��&������[%/&7���]���/8coԃ���}�ȃ�7I�w�VZ+��f9�rpBz�#d�c6$�w�����cDX�y�G�Vz[��lJhh/'��O
�[�^FS�C�l��zc6"�W�
τ�����N@Pϵ�ډ%Ų!F��h�����'`+��q�}@B��7Ib�*XaR�1��H��"�SY����[ �w�Ŗ����79/�|��!ۇ�J0��s�G��I�8�7pv k �\�ˬ����x�v�1z�mF���5
ɓ�<+��q#���q�+��ˮ_����� 32
�B�&��ٲ̚���Wc�[Ѳ�D�PR!�҇i2GNn��oPI��v{:pÈ*��z� �.e��h��]#�O�.Ň�ZH�����l��\��
�Ny�/�=���bVC,�I/bW�o���H<����������$e��6 #`��r+�zF	�ת�	B#�s��9�[�����A�Y�Ǝ�=�(_��Ǜ�O�4�I��"�Q`kΝU���w z2��L�(�b��HG��w�w�hŊ����0-I�
4����&�&3k��x�&��qn�&���R��%��wB4�(�p~��� �	ey+���U;�1��eKI���Rb��'�LV�V�o�H�E2Qi$HW>��K�@��p�P��a�b������=�}�� ���%�m:��y��(�H��D�� ���<�
���@6��G�S5e��7bk��y8֛ڇdgw��9�7�>OsA*J�"(�:�pZ���h5���QLG� ��7�1o�i/���D���řF�N��@���w��NQ��N%+�������X�%N�Ɵ�YC�螷�"�����t�.#�N%�y)ȺH	�X�:I��x�G�� {/'�;�����N3Q�Gg)����E�����l�	�s!��,���x��"��"�H��4 ��;��d۬�*�E��&�I�j\����E߭������T5o٣��P��h�kt�qE/�")���? >ÑF��pG�~z"��*r۫p:�����[���/E�v��'����|!̟P��0�F���Y8 2�:Lk���D~�Iy���8���g�T�A�fd3��@���8D2�����O
�T9/a;�u���W)�>V�t��:X���l-{7�AC���먶�7����)8^� :z�o��C��Ay=�ue�!�y�@��L
�U��}V���'�֗����q��j�*+���i��x������S|�f���=V���=�zJ�~,G���H���#�N����m(�I�,��5첕9�t�� />��C�<;T�ng��K�����	K�	�(�Y�����v��e��
$!]<�t0�k��;P��ЙTP`I�)��h��Y{CFBO�ٙ��)B^q>J�	�������d��s#�իO,�O�Ş���v�l���W��P*1��T�wWV�"rJ�'�R�6�`����)4�2��.C�c7��s\\����]�J��s�`ED�6�2c����p���y��n�ض�drR	J���v{��uF@���F�����:J�z�ܹ��M� �v����6�%��[66��~e���5u�ͬz2���ň���z��|�صy�!�$�f�4Td,-\Kj�J��t@�<8;b��15&��2l`����5R�J�|�j�k��9{��+|D�s�����@��8>�NU'�OW�^��C���f���
����o�+K`$������E&Bw��}��P��)o&��ޚ�^Or�k(���E�=��=�"�r�^S�I�q�Z�� �|w)Ff knr��g��-�F�(�Km~��g�X 
Ϥ�3yD�u����/�PnDCq{~��)�%���3�	DݳiC���NSi�,�'�qO+J�4�1��1-�G��m\�u��WE�|K���P[�2��*i�!z��w�u������ڥug���q�[��d��U���FnIZ�l�b�� ���A�D�}��u趌�`S	Ù����b���q��e&�;�^��N'ܾZ<�3�ΰ;�)k#�I�6�������M�6�E=�F�-4$��],��;ۨWS�Gv[��r�
3�m�ĉ�R����ǝqM��i#2tu����%�6�ze;܄��Y����2�-Q���T��������9Ҙ|5K��(!�A��-�/�W\��m�3���z�Ae,��7J?���V5�G�3�׈M-�+;�P���8-i�?SJ<eC�����3,H�
���8
~ ���%<0dM[�a�Rv�@T������ �qy���ȱ�]� �&>fa� IF� χ�چЎ�T	ُ*B� ��g�Ṗa�Q��rK6J���)�I4��[��JD-���i���!lfB���n�be��}���qG�o
�dW�X�#8I�i��!��4?�C@���1�w��ٺ�uR��K�1�Jj�]_�[�*�b
Uyj�㥶{Qt�+z�L}�`��S���"X*�b"���eL5���i;w?�U|��͈#�
�e���T�ځ�G�x?�dH��̽��7�'�d��v�<�#��^�qѶ��� �)����ۉj_^�6�+�/�/X�fG��Y�&�� �a����盬��Qz��1�`�J��_����)�����d�D������_�e���I5J�7��~4��[o�l%��l�,B����k�{Dz�B�8��fN�9�E@P�멧EQ�>��T������N��a�[fL�r�<<7th��<l�W�cF�X�4s�i��
��������%���kP��'�q\��:��:��2WZ*�'sDܵ�;IW|16�:�IHֲ�%�!�pDe��=�8@H�àZ�R:.<�d)�6J�	���5���.7�md��'@��,�}�
�a2�Qizׇ!����r��lO��X�"!�y6G��i�X�*�)�K���M�(��X�d���c�0L�[���})\�7����_޸����c�̧���[�C0_�Br.�Dr	�V*����9�5d���2q�S��2g�(|�Pq�xZ��Z1�1a�ֹ���=�Hc�_ [�2�h�/`!G\���̣-Y0�z����N����?��0���fvO��&oY�_���q����D	Ԟ��W�ҵ�t=��6~�S*Fw������`�2cCT,N�%�׭J���
��c��zG�����)�����Y7Gaˌ�Cָ �9������#XQh슷iyﺕ��,M/p3����Y�TCl>�Q�ə�����%ovY��@�!+,��K(�)��$v�*� ����U�͔�1�:ς�1_��m6.�R�K�+6�}��W�K������BK�s��������=Ь�=5tʖas�w$�%�$:��H�2�N�k"�<��NJ�V;��� ʤ�(�_�O�~�?����ÕLG�Y����M��l���h(�zLi;�@��p�ٖ�!2{ڶ>#N���K	mx#܏��f��*�۳O�L�g <�d��%���~����J�\�ώ����6��:��`�Fw9�>��?��OP~��hw<ū9LJF�wE"���; �GA��@�{;:S0�9��Y8
TpKl#.���;���4���9uV��]�GN����a�(�v��'��@���\%�A9��W	ge��1?I�Y��6�\�N:���m@:����M��������Q�d�F
��:y"N�~��S�li��Y�V8�EUBK�A¨Z/�4�J�Y��!!���� g��b��pF�#$���G������P��otb΄�ք��Bv��8?��+8X�O:�V��V�ᔣ�gl�:3T0�h����G�(���ؔ�~%%��roƁ��l݉٦7؏�����D��w�D�l�-w���� �G�ތS�WƝº�9�i����e���l%�����qTvH����M�o�NwA$�eF�5��T��qMd��n�f�M�����Tc�����[�<mΎPD�YT�B��$A�'˫:vQA�&N�F�<d���7�f6���avh�ÃQ$��	���(i�#ՊJˬ����T(i�CnJsd�h��O�p�Řu��+m�.	Gփ���B�!t��
Bo�C�����Ќ�o��� �:t	L��nLi�Ѻ�m��^b�'I�vp�������N��7�R�ɛ|SK'�.�Ig�4j�H�G���
��q"x<�7�5����I�s]!~�����Ay�2"c�-��|�\�%M+���o�����]�_���%��>-�H�T�o�OUR�����~�-륥�4�gp㻊��kl� .�80��@�W!�5s�K����΅�{��q�Q�����Q�c%p�Q����;�
��{	�N�����~N��S�M	g�B���"n�<�`f�@�HO�PY��f�t_�<���n]U�}�
������u���h�
���?�Z�U3�#�0Pi��,�<5c��r�ڤ���9��s�k�z˛Qr+�z"#P f4"����5J��C�E▃�k��zo�Ҵ���h��ۺx�4��	�$wo�M�E>���z��`(��R\j_��T�I��+�f:
��k	�V�͆��yE�y���b�H։tzOxV�.��r��!Z����Լ[�5k��w��[�FҼ����C�?<W�xjO�ޞ�t�L��5��"t4�B��kdJ��߫�;="W�K �����U��^Y���C�O�d,׋�O��&	w̘��}����&k>�H�D�r�܌�t���)ك�X��Nh�����1ԃy��8��k��}�%-�M�������L��*Vn�� �<D����g��-�|�f�r��en�t���zp6�;��Q���nu]f�㤩�_�é'����U'w�Z��X6�sSP�؂��# ������e{J����a�%>�-�G��Wc�L�!��G<M���l^K:���q���C@��ê�4�g��b��Xp#7���b�[��)��#���-i5O��\��EL���o6����V�s*�#WcRi��oa4���H��&��d��	GM��@���)�E����@���2F2���5�p �t��n��`�8���������ɘ��P�X�)�t�'x�y�����v�D�G�t@L��Oh�R8z�ɚ�@Ѕ��p R��/�3�n�?����߰�m#�HO��O�UN2k�,Β�^_�0>��̫�o2�`&0��L��bޗ\�׬߃�-Z>����R�Ttq� ؞&�U�6��$�!g�����Gw¥|r��)�F/#o�J�O��X�2K�B.�Ϝ��"������mB��f���pՃ���u��Іd#��S�'�����J"$79lڮ?�9b�I��%��8�a� z�xD�����4*��J~�*�8O5��n6n�z�	��a�~�&6�|�T�������`mT������}�%����8lLJ�
�e�].PU=����j��fNﭐ�w;7'�G�͸�w�V(l#�ݔ��:�~�y�K�sB�:'�Q��<c�3�~gN����P�T�f�����@�+�{)cFdQ�����<Y�kPƟO�:i��f���TȜ�?����h��ʣ1 �~<R���
r<��_�R��_���U"Na�f�6I9@̌�d.��w������6�`�Z��:�p��_pv�N���4X);�HW!F��l5��?D�a����$�[1���S���+�i��n�����{���c�6�o$�c�ZkL �6��f��n�1e��*q��U4S����ZW��s����ltd��J_�(�����r��NI*{��cZ�nEC��(ڂ��oy��WF?�"�k��:ȪR��`��6���!/�)�uw����#��MJ0(ʹJ:O��,QD�n�>Z��˲p�
���N�Z�G�R�����"��a�:��f4wB��Jp�ɠS]�� �\�bլ��$L7;<�f����g6��OJ$��:�pJ2k4�7����4n��������U�p�6Ԑ�C��k�5����;ۍ���GH�/<�3�9n�� Aa�;>o"�}����v�Cr�Jm�\υ��2�VAv�>���v�0���Y�;+���Cs�/�ZU\	Y�@PW$ٱῃ�W�K�y��S�j��q����j�"�lX'8O@��?���S���ܪ_�%Az%�r���w7=�g��Y&�����)	�[��'�9��叿'v"��A�)����YH�*};13'6�ڪy9RA&�\`"Mۂ{Ck�}�F묁l+��|r�hܢS�gbS/v{��{��<��2U���>Ұ�h.�'�Emo \#�#����e�zX��=k�8�-�hwٞV����}ݳO-'���d�&t�g8�~s�ǀ|F���dF�ʮ8a���x�@���ze��y���<)��%���t`��h0��o�q��&ʉ`�_B��e����<p.��MD�c��YCJBb�T� {N�� e�d�3��\�t�[��k����aw{�'���"���ƕ�s�F��|�H8cH� �mV3o �2����1-,���i�n	諾=R}��&ǐ{�Y��v_�U����;����V���O��U��m���śz�c�{���E+u����"V}�DzBb�	���U'��[�,p�!�pr��X�T��.&���8��l������Eic���4NK½x�2�?�vLni�<�4>d�N�ꞝ��{��|Q�2��{t��v�[lFw<�e\f��@�V�� ���!��#��Sp����#S���%�T��J�+gHCi�s��.�gv�u�ճb��!K�P��2	
��:܃t�P<UP׶57�w�pP�8��a�l¿a`�������t��w]�}�����I�ڱ¢�`�޲OKI}�[l�T�\qM���ۚ4�z�p��M�U�.&����-��}�����@0AD��c��%��)w�\뎞�Œ�/"dP@�M������0J4`	�������A�Ff�tX�r|���\c-�������!�( q|��Ra�K�Cnj�O���c��,J���+�͟E�ż�����:���0��bă�)�ױK-�g$OO��H��p����m��h��J�vU�4&r�U���<���^V_�OAi�[;����2%;���4��2��J4�g�nǖ�h�K�&�˥b��W�dsxn5]�DϰP�
�|(X���@��E��]�y�(����6���nĈ1���s<�4kF��Җ�f�����,�@�9��z��U�Ť��mz;!ܢDfux��3���J!���8����]tllA<�n{D�����E J�]K�JZg��=��&{��q�7!K)>�������7�<T�éf��R�m-t��)����[�2=����qr�3��o�q� ������J �F�1m�if�)H�6n�R���h�/O��1�F�AK*t������fC%���w7l
�724r��p=��6wz�A����p":�4����������/��YLm�)����iƜ�n�_q�R���$&ڂ\Gk�罼Sc{�=9~�F���IT*�^&hЕ�� Ȟ߻^-�z��b&8���ܳ@�1�j�ϓ��l�����{`ɉ�oȒ������"�i+�����m����"%���(�̃o�V#c7�/2��7�&}x���sf�q��%����#c�=/�}D����t9�t�N?I�5�f8Nj�;��c��G�*�v�`�k]�����g_2w�&��bDr>a� @��r��ғ&9Ͽ_�U4"����୞u�Sf8����JY�xf��}�?�h�:tT��^�?���Sj���ePH��d��d������G[^�0kE��$RO$�(0.�T���9�5�G ��>�&/�1-'5~b~,j?P��0_237E��DJ���d���J��p�������[�"����0��Oܜ�ob��`�H(8�B��:<ۦh���;�k�5u�<��ݠ������:�'M�~_g�w�!WH�%ǣ��&p8\���N���qf]�f+u��f�u�fr���9.�V�h��]�R����
������I'��HrHGs7-hܒ����+ڰ���c����}���[��aQ	��_�P�"�z8Z��S۔���.)���t�3��{�n�C냇j 28�lܥ�a��n���x�!�J��ݩ�bz�v����d��*��%�07�7ǈ��%��WjG\�bqHg���ɛ?���{�4��T�{U̧�62��^2��;�<�l��:?��L�=I������T�JDjl�^"��Xɚ��hYW�Bd��4�&�%���a�����k�I{��w�.eW,]�����R�������@2,V��FD]�G��V���M�yD4O=�d��,3���		�6P��V^�R�q��@�UfY<J9~�O,�0�� .�|
e�J�y���鉇H��R�ыm}�<���QA[5o�j���i�1,I��:���a�R�֝�1=<�'�#h�S�pf��ۨ��+�MF3Ud8�C߭��[�9��[��t��[5)�cx��y�㢆H�Db�Ԏ��W^1"*}b4�A��o��J��F���.�w�3���r�ha��%K�v_�|�nUBT�Ԉa��4��!�V�u==�zϬM.�H���;Z!���J��C�nW�X1��LR��D��� ���zs}Q��Y �-4Y��4Oc���Q�� q>`S��0�/�K%'0i)����ߓ�e�L)����i&p8Bs��h��m�w�k��-�.ru2G���fʗJ ��Ԟ#W�Q��[2���LGPt���wS#4�O�����oi���C��$��
�:�d�#��'j#����y�9.��%V�>� �������
��|oT��x�*[%�eN�[!�mī�߻-?���h��%�d\�vOd�@����'�"���r".z�*�S*�>�qIxӣ�d�5��;��m���Fx�1�Wn�;�4����ܚ��i�M뀗�X�;���._��Q���_�3��4��f�
v�����\.�UA,��~�:����ࡐSN�t��Q*�R{w���D$_��ɒ�ب�,�	? 6�_f��]�J��	�7�yP��Ő9�P������^E�v�j�VJ��)���1���G6�Zz�Vއ>��|n슇��5[@ǋ־�eN���𾏇d�
x'�˦��p��]���<�H1$��ջLp��n_���Y�q�4��H-�����V-�J4��^Q�j��E����LOdŇ�������{R�vX2�.���m0I�kj.����]U�.4�&<�MOHKtPtK�m.�T.Ѧ�K,脿}���'0ԸA_x��,��Z@�8$�������Td�`��$iV�t�+�#l.�m��IU�w�{:�/~[�l|4�;�س�B0�7oY���eq͆��!�h���h
8�ՙ����^y��o��Wխ��|��K�g����ǔ��)�.�4��lv�k��W�k-���ݽ�J��f�:P���$��<>P��4��:�����0.�CK�z��I'o[�9�����
̅r%�>����:!A�Ԇ}w�&�G�=K76��X.��t�zt�;V�� 
 �v��.5����ZF^7t�P�O�x��M5�+HH�ڭ�4���z}��
�"�(`�����2F��Y��8߃����G��ǝL��tj���0-��b%@�c��PѸ��X_�����L)0Fw|]�l��!����k �WE����^er5 	 q��>
��� ���5�y���x�"����-�������zB0�<s���k��4f�lO�a�rW*e��H����`��M�����P]4G�J��kJ�vm)l��7!m���������U���O��d�/ۣg/�B�����w��.������M2��>�
�|�Ev��R?����j>��1Saݙ�H�kO�G�$O���]��z|6  �E��􎖍��{�������ݪ���鰔����̍����z-�f�H��dYȥ��V����Hq�L���G$���uq�Ӥ�����k�.�Ľ���0\8���b8%��}lINi_�\�|���<����x��ÓD�KW���/D"#�s�G���2p�-�gp�Ŧo {S�2B��_��4��s�Pߔ����k=�x��+���̨ɹ�[=����㢥�DW�%��S�6�H�WsP����s��O%��V��!թ@�[��7�%����rl�:"= eJK�!7��ig��}���jQ��ݞ����'��T0\Ո�Nǫ�=�_$u�H��ʖ������j�Q�+YӬ�G�2��+�x��h΅��4N+U�� jƳ�h%lzM���,�a����)?;��9{~�vA��[�2���o,2�+��x~�0���*��q���M���?4|T��bew(uɞ0/�~�&�K�������wH9�m����L#f�����"1J.��	C%����)��e��\<c�s֜S��5;.V
�RE�W@ ݹ�r�M�ed��0�ֈ��9,>9o�5��⊮�s��_\.z��+���w(�#�(�w�`z>�M�?��9��&#h%�4������=�)<��e�GΡ����B���#A>�Sy�v#)�#���|(�;��.�g'������v�H���Lz��_Rl�S���Ȣ{�\~�' &l���NY'=/j�5��/sa�{����[�̈́��q3a�E�#����#ީ���?1�3�;�U3�b�Q�]��
Ic�|����k�r��� � �e
2,JZ�\�8��l ���1�	sMXp�l3[}m}��`�X�?�c��"ȅ�cL:#���6�RI7���e�Cd�KNl��)�gw*e��4��$%��g���3���*M/��jz05)~���iV����h���mGG�0��#�����ç	3?W1�R���� �d�v �0��^�E���^�*y���>��t_[B��Jv�lL?�h��Y&@K0l捯��[��K�ś�֎�����#<8�IJ|�~(2����F�/��4g�ӿ��K��ܭ�A�GO9*�^�h�ի��T�Yc{��#K
dO�?�������LE�qWo nF���2��2�Kț�ξ��m�Cmۗ�FN,t�ݛ�b �|�Xr
��՞	i�Sw�Dǳ����
QF	N8��-��ۜt��^�WM����h�e�e�~��� K��xMδ|���.'�9H	��� J���߫#� �>N�GB�7�B�b	w/`wc>�nE��?�����:^I���m��Q�#��}��>u��ű��˿��U"�"���[��d������~�D��Z����W>���Өm�_̼�B��_~�{���$�@�J���GŲ�5Μź�O�WA��eLY[�jOg�Ş��+�3��}�@_����&x��+�P~A1d;�IƳ�
wWj��$s8,f!J{6ܽ��]9�O�5���n�a�	��2UM2�^=�$���y#���N��v��_�{$�1��'f��M]�d��-8�p���F�]אK���l�����gc&����ʄ�ݚ�����΄!��CM�����(ɛ��܀�Y�C�]�:���#`��.�Q|�[إ^�!5��dQ���`|NSt�Q��,����7l�ozỳ�n4?(R���v���n|���.�Ҏ�2�L�܄q��;/�aG��O��HK��Xk�]*�kϓiV�.�I�Ò��X���~�������up\(T��(W�G��W�L)�� �#Yr�E�~WZcDs:.��]��Ўx�x��.O��P�ߪb�b<�|��@�b��NBF(�c���+��qej�і �t����1q�q>��R�)G�^�˺x��v.�� 
Y�=��0C~�5�	pm{��9�������(a�u;��mL���(㽭R�8_���^d
(1	%=��{"5"� �������-���cd}�ƒ�>�9�U�ɋ����!-=-`h��n��Tܖ�+���9'���^]':��]���*@rvp'�6�7�`{��b�&���yV}J�
T��F�aN\�j�b��e�1���:�R�cw���hB�A�Q�ظ�z�������]� e���]�Z�"�;kqm8d��Ks�	N�3_�~#	 �FĖz��N���v��A8�����|p��B��'<6�����/|�u���Oޣ8�s6�-��d�P3���!��$�a�?�o{^S�@���:��ͪȫ�$]0�Jl���ꠏ�h����d���;�T6�S�[�L�N&j�<��F1�]Z�p�ʾ)�cD�l��wԤLR�m�>��'����a��kqh<=ǽ�nV�ڳP9�^�a7��&��QsU�d

3_V�%��?�8��~.�J&}ϣc����EV�P\OI�O�z�b��q6�� )�(G=��m"U!$
e=���$lh >3[|h����Q�*� �$�Z����yY^���e`�L��Mu��.G�8��^Ku�o�J�U�Sl��J� $7���U'�U1��N�� 7��~v:���{UuP���b�j(��??皪b��_X`��Â-\C߻1�'��Cͽ��	/!�s,�5��F�=ŷ�_.�xI凵T�s��
N/Cq�LE��	z��R�QT��f��.V�����Lx|��~��F׺�/5|0͵�t��.��z*�Ҳ ���(��C�1pQ�Y�!f�1����'����t����j�'TA��M�_nw��}+�;ӝ��Z�!�R������q�H���
Q.�d�K!W�9�hO�R��&+��l�c���ƥ�SA,�[�~ s�.˝O�A����s�i���s!��*].�����k�XN7G�"+\g�1_����><K24մN��Wb�ɢ�],x�\�?`kXΝ�Hp�4�;t�ne�q9�6#�"��	~zY��:v<���?�����,�=Bg���{lj�w�uZ�)��s��gU�r�;ј���3��(~+��m��LK�"�r\Δl� �6�]&x��)��)�ZS���xv`�r�m�S-E�SE�/O��0с�����5s�h� ��&�Jo�g�ϔ:j���u��Aٕ�H��T%��_��;8Tl_��;��w.�,[�uSY0�HP.��4����*Ư��g�7vn�^�;�}2��$�^��-D�V���by�y.�����ǡu'�/��15��\�{ԏsՉ�(�C�u!��R�gёI��<��^��hh/𨓕sa0a!�ѓD�Ad��T��Ty'W���n1#p-9��,��}[���~܁R	�W��(�|HnBE	N��Y�Uן���8H�*�z ��7��蜇0L�azX��2S�"1� V��(	eC�[�%q�������������`�\p��S�I�A���B�uӷ#~���Fr*�O��$w`�f�0[ކ'̌�z�dz��:�zrM�	+o�6��!�	g7��ԉp�^c�#�{E�k�g�������M��[�q�y��٨�3c��	��@c!� ~�Ⱦ,�r?���Zt���Yz'���&��<;��K2UwĦ%U˵?r�t��ܴN�Pٕ��|�pY�u��L�"�Bs���dE��ۣd�Q� �G튒l6���^��W������������;����R��E�N�����=W�n�(��Z2����K�ҡ�����3HƕP���&OI)���z����J;�o*,՞F��ݾ�щK��� '�Χ��	�o��r�&/�&?³24;��s,�˄���ⱂ7����뱮8�D�>(i��-�|(�r�c�xW���J�{�}|�5�yǮ�����]j�ͨc��^�����7����+t���^�I
�^B��'.��h�"M����]�;��(V�%�׉.$ؖ���I(Mp�0u��v�}��K+䊸 (��������SL6�٥j�>�O���q�@)BV����b
SK:<�5��> ��ʾ�l&�;jƟ(u,�/�4/�����b{ce��GťwʈEV*��� �
�8 �g���l�[�r�tAL��/
4��I�ߵ��r�s;<.�&=��D=Z��D܊�qc��;���6��;�7y��x�N�u:�@�o1�Z�ŋ����<l2�oU6�ⷸ�5 �)6�S�f�n����Ӧv�� Ϣo�/�ߎ�`��u�R�܎%�/�OnD��~-ߜ],qٟ��4�t�
�-E��&C���M�C��匜�I<R�0�u�ɁH8���%��si`������'�`*�*	�ſ\�~���ɥ3�����O�4o�+�K�G��
��`E�#�!O1������+ֶ�*>AB�e�(l�6
�Q�
�fɂ=�>7�{=�dpu���eH�F���m�i�DBq"TF���������f4%�I�"F�P�����^�����+���8oRF�К�q��iB��𢔴�D%�*���&fВNV2HM͛�1���5����F���	��1��T����O�lKx�|*V��k5�{��s�MNcݐ�/�P�r
+����T����bb��t�����ƀ{����]uӓ]�7�1�\c�	��M]�]3��S`	f�]�E��\$�@��lp���X�!ǁ������Bˉ�aȱ���u_��Q���v�J��[)ipn�{��N8�%$��D�uLv�X�4��MF���80Xb��ș][J���O�7"0�D���ǑsǓ�Ż��_���E�u�ޠ�Rw���h�ۍ���Z�d�$A�oL/~.�e6U�&g�r���DW�Q���}�Xe��J�~�R}�m �AӇ�k�8�C�#�ˆ(tP��$�m�4 <1A{�)I�A���h��OXI�{Pу�?E\1o���I6��h�Z��$<V��F$"�4���!�8����4�\�H y�Y � ]$f'7CP��P�R_AhH�	9� E��E��4͇�X�ߑ��R�������Ã��!V�C�p[�-ʫ͍ m{���%ޙ�y���/������_���"�.���6L}}Na��@�\�2��q���.9B���ߝ;4�A�k�k�_�g)y�f�,�.�� �U2��+v���� g��i�Y���S�rF ������)�ߢwf�y��s���ˑGu��1�p��i�_����}�W�g.~�~��(�\NH��woH�2�R�ݙ\U��`�ј񶓡X�gP�ܕ��_�����S)J;%����oJ�n7&9�26	�^�p��M�m�b��<�_���K�M^=�Ю�(�����O��2�/���Iv����Ch�`�&�/ő<�?�:�Fɛ��oS;�FR�ݩ?y��:A;e������gz���>7��ǉ��Y�$�p�H8�u>��<�nM��6�`�:�,I��L��)r��w�4r�P_�/o�s,#���Zi~s�@5�U�,$u#"�{�X�e���&EMB$"S��� �a/��삥�|�a��E���B�""� ��!���<��-�|�XX�}�QJ]�
�!���(�2�u�_ceYqR�5`�[���m��k�v��.n�D��DJ��� ��֩���6۲�3�cw9�-pD�*�pAT�<��<>q@��<�b���i+$�2���!����5�Sԅ��f9_�`��B����Jw_�/��
{왜�6=�;\�y�*y~�,���{L���i���S������[�����T]Î�w�]�)w0���$�����k�y��)������\��*@X砗+> ݏ�R�;�C��S�<%J܊�"
���^^`�|Quw7zm�"���E�	�ᢾ]����m�?�r��H�)]�D��z�3�)��Q;;̱�4ͨ�ӗ�2���D�o!�s����~�7E�^S��Qw%'���R��Ĳ�F�px<\Ը�O���fb��,P���g����M�m���h��q5�Ao\a*�A�G�e󖊰�j��K���<`��*���(m�C�gTR��0�D�c�T��I�Y�l��De���}�Z��	���l�`f��¦�^;㏛�Xr��r��U��&�_�U6^��y�j���8W�X\��C���T��s]Q���2\��"WT��e��<z��PK
"�������Y��i}Xw�<Ě�Nߒ��^�� �8W�%ɗI�K��9��ik^� �'sZ�8n�;���S[�_$��`7��E�<m��	i̼dr��H��f�N:�����U���aڀW�(<�bf�$o��\:�����-�J�w�vyC�:Cj�����ʘ|�ؖ���"���iҖ%%W�`���:d�~���G]&��K(+��0i̩H7�+.�E�a����9Y(�6>�T4�t�e����jo�)�޷ތ4���b:��|E�:{�A��ք����3�
��;�A�f��5Z��h-��"d(P�3�>*ZO�M����6Ѥ"�a�؛z3�umw��{~4:���!~s�
*�\�q��C��%���y�Y["�l]b��@�^�)'A�)Ɂ��%w[������%Ïf��5�:fTk������	
u��9�}�&]#C RBg��B�ك�"�c;1�N�@�RC4�Vcc��AtN�գf(!P���y#L��/{�����0�ˉ�L�����M���.+.5���VNd����i=y`6�o(���JTln����q�l�N�*�M�X����bG���l�Vo'?�]-�xr��1#�<�K���py�>1�PsXz����IZ�Y �r̓5��t~�U��0�3#������r� ���ؓe�;�v�6G9�Y=��������i���C�����ƞcئ�Q~ˇæ&���!d,��r��S�������l����p���dW�N�a)ѶR}d~��.�o`��Eܾb�7�j.l���H��@���=$�k�rHo���oO�Rs$�U`�L:�&L�
l+��0�^qO9���ekA��g��L5����ՠ�
�25&���v�&V�� z:Ԣ���|F�٘7��[�
�l�{9���}6H�9��<x�z~]�9}X!ҪW����A��yc���0��O�P|,��"@�lk�t�f|��Lᯣ�cǑrGu� Q�^��m�{R�"�qY߈JU2׍@�P7��{<����cUe��PX%K�խ�e�K0ʬ-�hDW���%��^d��86�ڑR�)m������Fw��`���눜�Af���+>Q�h��I�CKC��E��y���S+P�������x]�ʝ�ӧ�}+kء����|%ќ�Ƥ��v�cO���)X�R�m����v+쇴7Z�i7(�
az߻���aZ�J~�)]�@�۱�e�L��V�RCDn��\O`8���7<�]��txm��C�{�����mlL��#��l~�����`�kg@C�v�xqբd����Xg�P"F�4d�z}�At�@�w�EE~���ΘWХ��!<�#�pEN_e'1���r;pt ��
ai��w�&�=u;�sW�y~$��й��B��Y&)��i��l2����E,Pi.�Z)K�-��o;ٛ����Eo���ܪ�Z����an[^�É��V�D�f�ٕ�j��	�K[�g)e��XѢF��%�ўD~Oc���� �Ϛ�ګ[������\��W�򓱏���%QF�{��h�A��w>���"�,i���vZY�>�le�OXR�3�����G c�Q��1`4�c�i�,*`"�JɏƥA�s�wY;�"��K��.f��~5cL��=]~�]v��QL��őnU(�2a	s5�f,�i��;YX�+���BA�������-s��S/ӝz�(��y�0����ȇ �y�alb�d�t!���0m�,^�-��7��{�V�/���b���$�	��%+�ӻ����U����-�vG`=�re�\<��)��q\����#�����R$:��;�j4K[ܫBG_Hb���}d��c�
@����gtdG�оm�zd3��%�����r�@����[xF7Ȉ�x���t3�|I�����}��|��R�pUk�_�� ʗ��FI�R6��_��˴�{�C����߻	���7�R�lvEzS��h���cy�;<8����Z�".@��uS�l��Q��^fG	�y�e�3�X���A>PL@s%@�+ V�G��8"}�:[�8���i\��=��J=]��Ԁ��a�?()q��@�D�g����D���!�Sj�����7#,��>?���AD���P�|�z2Vӣ����1ܳF�rP� ���1������y*�6|�x�EY�PÖ��C"݉�U�x܎�G���bMD��^)��@1�����d�v),SEkٰd�Y�X�>y1���_�����q��J��
"B��{ŰV��8J�p[���u	�(���S�|:Y�3����(6��Q�,�g�$7�mv]'�L8a�D۱(
���_�A4D[��=�ɻ��Jd�Ҏ?(��g�"��wTGF	�#ތ�F�Ъk�㒺pva"L���r*��v��K�(�@&�����`�ߜ�1H�v �.�q��]��a}$D���8*b���?Z���>��_���dp�UMS��x�[�SH2:��I>��:�(��ػ�h�����Q�,9�]��컄�/�xX��f�SlQmR�0�j{a���;w�)�P_�*2�Dw����26��	���kE���y%�sd��Jx�I���'��+C�u�5L��YI볁�[���q����T��?�Ѭ���K�[LZf�����,�R5�+u��#� �ǵ�Z��� FO`8�̪�ˬ����.C>�>���Z��B�NhQ.���"��x떂x�MU��(֞��d	����}�1�H���H_��JK�P�*������UO�c��K!�G�E����pMcs��2s��:4�є�-�B�__�՟�]e�t��R����.a
X���
>�]�k�U�pZ-cy��(��A���sx<#8#�n���HKN�(��2�n���0"�'K�>|�'��L�5Ԭ�h�3}YC_�%O��r�w=������U�	,iZ�)�"��0�9'Jt�m'���M#02�1����x���^X�ŗC3�i�Н4h�מv�ߙM�2{�h�w`�P��U�Arz�d0+8�F�A�w7c�4pQ��ԥ>��2��OgӼFϞ�c�M\�����$��~�݄�K�g�������]<�Hl�1�W%��7�����D�jXY1�=��Y�)|��RX�#m�4�:�����<�/��7�����Z�T��q)�	R��U
�Xʱ/��K�)v��<O���ҬϮ�ښ�Beڞb=�f��]�q�e��"�1��:�(	 )bI�U�h�Yp��q�R��,`����,����O��_�c����[Qkx�I��Y��,KR�8]|�W��������A�LR90}��I��S��ݡ�}��ꆤ״�H����VMd�%�&s
�W�_=0܏�j(?��z��4%��n���p���~O�����}4I|ɀ�����FL-PrFU�k�fI��}�p��f�`o��s��� ���=A��a�3���x�<�����ĺ:Tt%3�.�v[0������&%�0CV�Kg~�OF\U�%���JmeGE�WG�h�n8o�A<��վ���EDӝ�s�7�o��V�P:^J;�P� c�����)[��h9\�Q�|@��c'�K�����]�^�#X�J��TH������Q�����a����T�����iP�=��T�Lh`�e{�E�*�Y����l|凷,�'�^K�ᘯ&�������Q�+U�ˌ���q����Ю4JA��Y�!k��f��������''1v��]�V�`��ϿFr��i�Su�-v?��w_�����"��ƬŅ�A.0�G��0]q~�S��ȟ�P�
�����k�jX�e�oq���zZ�f{q��w� ��Aٌ2�9�=��^������f?�y��¾�s;�i�1�m^�٣w�������������#��4����5d["�[�QX�ܲH̈�4Y�4Bm\���kP2Q���;$�p��g�ʺB4������р~G�Q�N� 7�%�F9�A�U`J���S)���
�^��~4٨�դ���Z�b�e#"�^���B��nNX�e�$H:�Rw#��9��ˀѐ�;�愱�0 g\���2-b����l��`���	�����1"�5K�����}�������&�o��Eʏ�nf�N�JB������e�E�"�se>?�u`~�U�D�x4��N;�!A�@Wa B9���.�+��/��s�z���1�k��
��7�t+��T�[�;��0��bc�Y' ���H9\��i�zų|�r�K�?k�������(VT�jO}ue���қ�����aޤ�M�Pٌ�l�|JY^.0sj�Xo)"�[��pX�y�~I	�#�to͎�\�-+��J��%��_� "x��(0,����)��H,�χ@�[F�O���^�{�%�{�H��LybY���w���aɍ@���Q����!=�A���_��(�N��Jq�}��X�j�����j�6�����_�0oJD�/j��;�i�X��	��nJ�Au-����K���}[���� ��zC�n�S�g�'z�q=�ą�P��$�(/��,J!�i�&,Ihe�*�Α�@vFp�C��[�Ӳ�
�die��ƽ��$����?o/I�K�d|�%R�t۫GX�yџ��|.��\y8W��$���-ܦ.8��8��2���e�H�Q����W��6� �D��s�Ǝ_T��nڃI�?��k�|h����u��(�r?�N}��Ǆ(k�K���"�%2�:�-,��#U�a����x������b�>O��YN�����@a��ᰛ�{
X�+���s릡δxw�]������x�J��mϗ�%�4��5Q������P��� �ζ���*�B��`�;u�Jxz��	؋99�H@���s>���|�����z	��z��1�sl���>y�pIdޕ�ƕ��~�'u����j�&�e�w�+��*���9��PH�V�̆ꃪ�?�ӰqX��p�Z!_0��^ أ"tP��E<=1��#��4W"�u�@P�&5���c����T�#+���p�.�JW\/:����j��/����*v;C\�/���7BO����f������+��D�4�L�!ي�K�Ʌ���۪�Wݨ�oB�28[y!T�/��SBy�*E��N�5���]R�F���s��4?At�`R�ls]T�'�j��ބq7~��ao��&J�*?o�m�z�W�\E�=�J�|Ɓ�\r�;��D]�l1���.������v���� 	�o�d��U�W5����x��u�2���t�q^�1��߳�{,���HN�sr>|��CvԶK�>��\g����0�f^.�(h�^M��U!`A�Ćy%,#�gfy�+��5��Aع�.@�K�ɉ|@��"���vp��W�H���0BNҝ��Vx+	��ó@�4Z��b�U�A�2� 8�6 �s�,A�Ax�9VӾ�׿��R:Mq�;Gmc[ܶjX�L�ƻM��w1m�_i�v���H���s���zj�C�����U�����9���Gŏ�t��!cc<@�*��!*@B�uo��!`��g%d�X�z���;�a�����+d�5�3ia�M[�;D�Ղr4 y���Px�X���!e�n\$���ߘY�	ɭ.N��u(mAr�����q���˸1MoY9�~s=�����f�b^�k��P��5�T�k�V���"P#��@_~Ͻ�'��a�J0Y=�����9�'pg�D�45A�M��'�3QK 5��z(3X��+�Z�!��|LI�F�)��gU�V���e�ie;�G~Ͽ�����H����f 	Z�N�(Å��C���䤧��:ll"M#�^:�둯�@�|���Q�
�z����]N^��fDx}�Zܪ�P��h��DF|wߊ�DV؜��Z�������	;bU+��noGi��Sf��9^r��_ ��/��T2���q�'����o�_̷���)�;����Z҅K��v�.�UgΠxn��컱�2�5�z2��8�{�<�F�{�ɇ�*�|O(�2�zu��� t�|l�_�
Y�&�'�Bˆ����^�g_�Z����#R�K�v���
H�+��.9_�Bb�n8t���J`'9� ��Q]+W��e����|����z�f|OWl]X���I��M�7#��������^.���ֻ�'{ѣ�(�.�q^�{�K�J��4_i1$w��(�m��B�^.��R���5��^[��ت�U���\�F��U�w���}�r�H}ibRjӾ��M�7uk���ֹZI7������'W�&o�o崑�����?�RӬ-��s�����OR�M��צs�����#��?���3�b�]+�BOl����BK7vc�a:��5�~��>j?R>@C?�p� !��B�`N$lz�7xk&��K񆳺Mr8ݙ��Zn�$"~Ƨd�SK,8ׁ�8n���)Ѳ���f������"���p�����7#|H�u&S�X���|˜��ǷƆ|���?���w�c����Z;E��
Q��(1��&�$����m��<��;�WS��YW�/��8��ƸZ�����OX�G�ٍ0m�@b)i�X��mfK���ե7�:�y�����%���i*�c���s��v�"��
I�����l>��(!o�b�1�O�����������/��-V-߰ڗ5a���ӊ�.5����l���'wpͧ�����٫���#i � t`��~a-�'Y�t���m
�(�m�'XuS3��dɧ*=��5��c����2s�ؒR�}�1�G�Mނ�]%��B�%У2Ͱ+wjnnJ�xX���]b<u�iB'�O�����[�r͸�b��fr�;ퟦ�h�i�g�����|���)4}'��4�=j��@~��w��kb~c�\9���bvʐW��A��L��Fv�e	ٮ=?���_;n�~ۗ2��6ì]��Zrμ��ZQ*�qb�bҘؕ�K���e���z6&��&G��Q';��Zf�A������惉'\!h'a�-�V�W���oD 2,��iVA�[��	)B_��,A�:W���tI�!��]�TxAS3�Qdny���-�����Hb "0�û� CP����W'�
������Ȟ�E~X��tp
��9s�.W��J�F�ۚ�������F���Km�܊Q���'o:����wqX�mG�R����آ�]�`'�pi`2A�2�_S�4��Hr��\��Y&u�/$5� @�7��_[8+��#����~����G�$6�m�?��ql��� D��ȹ����f�)A��B+��Sta�PO��Hp����H�pYN]_��
/�m����X"���4p�q�C9H�	�V���ߞh��)q�bBГ�I���A,�ȇ.}��ߝF�D.�A��J�ಌ`*��-�$��X�>TR�����I|�&J<Ï�;�qs��Cx�A�|d��^�]�LWR$�=|��>���<���� ��9�K���W�bi��:wXڿ�/��P��y��K�#����Me��a����S�"��᩶����y�-��l���+/-��3?�w����z�^X�*>NM��3r�)����U�%��D�/�=�~�̙�؀�*�˪�ml�����rj�Y����r�l/��/ʒ�w��[���C{g%�l�������Y$n6_t�Ys#:�a�$��u��m@w�'/�m�4�ڱ��ˎ`��)��U�b�'G�1T�y�U�e�~�������+���;�����^����D�w@� cy�4����(V��;�@W���e8GK�����"t��➅���39Sd�*��g��Nuc"��Zr��df��z�<�9v5�	�������?��x[���R�ţ��zd���"��`ߤJ�%���;G�VPی�%զ���C�a��v5H�Ǜ�mj­r�d��ީ80�h��n���-<�[o��/e��V�4�Y�g=m��	喟�O����])�{�z{d�A��j."h��`�C�_�I��e&�E�f5n�n��*}���v�bLo��]B�EV�x����/�\� �C�����Z̿�	󋩈r�A~{Snd3g�5��B\�W�W�/�ӎUD�n�y�bQ�����G�s����[j�=U��F�dd�8f�^�����S_{���%��H_����(2E�"�q�Nj���f/p�ӺX��=�Ã�C��\xP��,��\�����C�F�UL^ej�)J��Gq�����ac�䉡�l��!���i*�(j�Mx\���u.�%��<n�g5Id3~��j2��''i9+����!��D���}H��|�,��G]�b�NB�2^=Z��?V����g�f�V�}������K΀����?���Y�|�k���d)^Pc[p���~��)��D�}k�L�g�+՛6�f$�P�ݎۂ�U��kQW��t$��P�s��FT��"�\���q�'ԙ{���t�ܔ����k:��ۚjG���z�J���'W<�Ґ���{z<4cE'�QSLJ����������qp��d=������w~%7�0�a��ڙhw_n���j�qy^�C4����@7�C�f��2��i�H^Ea����Z����,S����`T\��
�3�_OL_{Ȱ�Y������v�$R؃P�]a&��3�{K��Q�OQ�^m�7�� A:��Ұ�*�|=�uEu��1���7�io��}H����Ng�O�LXf�RM��ӊ?s!T�>�����2���Z��h��z������v���R^	���{��av���I�[�B��g��&�,�|}��:

� �霳ުi	���pqA-�o�o;�a��F��8�+��v�C��f*��O�,��8�&/���@�`ҙ��	�ht����9nS�aY��������5fAL����� `c��,�?����1&�Z�$�"����i�������A^��~�=$_EyiLU��_P��_�#͊+�f`5�A�<;l���F{T�$�����g?W[��"�Wf<a)qB�5�2;v�6��{ayN�_W8<�\ �j�M��"��e��.�*��Sڹ%jC�KG�)������VMj<)&�Ȗ��x�&�V�����mF����3�NBG�/�o��"�":�! �P�T��@<��aa�S?�I�|y�H�6a�QK�ߣ��텙�A���XM0N��~�0f\f��۰C�F�0��r�SWcnK7���@��),H� 5�[]�Z�l*y�)�V��H�r����|/z؆���;Z��j��RE���!R%	�}M�������.���058d����i�q�7�w����G7>�-�u��R�y$�L�$��BJ9�?
	���Z����0�%?��,R�ه�g`ęi4ѣ�W8�t�Γ�$�7�wEg�tr�0f�<���U_ݬ�1���m�<q2ؙOq=w�0�G�u{��p��(�wO&@���W�ֳ�Ik��8��"�Z�V��`���v�}�F�
�
-m��B�!t�0��=���X�� ϙ���:�:�w���٢a�J�T��X�>B��L�{�����1w�D5S����f�K�ŀ�u����`��������dN�$�J�&��y��12�3�U����v��~�������r1DT��1��i>H��(7�|W�mmU��G���";@EӨ6��'�h�uWDI ДN<�����r���@��|Zn�`���u�m���w$ ��� S�):�5���c(�"{Dʕ�:�#���*�Z�P�|��am�%��qi��c �~G��^�t��O�a�Z�W�8���!G���G9���c>G�0��G���L��=�W6*	/�;8�2ҳ�|F�<�Bs'����u<��V8W�l�����Y���ic���\���V�1�g�[!�@D"�#��FhN����{p��Wj�,j��:Eλc�<b䆩�!�y������ޱ���JC�)����j���AG!��aH������R�g�Դ���
�l��ݪ{�q*p}��B�����
;����k�|��e���������6e�l�>��Vh�wgq좜Y햆N���ח{ׅ�墛��
3
���ٮ����om�a�X�͛�>)#U&]� v(3R�U���"PQ̨$�����7��n��6���D߆zsi�7�V[Y��N�<��8�At��e�g/Z�$��ȉ�JA�(�C	��J�e�D)�E�S=SR� �Q�J�̓���:�Y�HȄ �3�� �Q򈗪�ԅҙ9�����ωp�:����pB�W���%���!���v[�!�K8	W��!��så=}W���my�=�-i�0����&ۂ�UM��[�U$v�]mn��"�詚{�-]��.�C�Ŝ�k�T�����wH�h�%�ĝ"&y&��PLW?��,x ɺf~�yZ	E�7��@?�N�m����� ?�!�Q7ezU�ǈݛ�B��2���Ϩ�W]��5����\�K�jz�Jl��]<z5PQM5��W�8�7*��kT�;�=���rj���}L�u�z������Z�`�gfI�b���ٓ��L��z�3�
�5�k#�[:L�Z6����;��l�`iz<�� v�ڔ���$q&|0�I���J�����ٜ�͇������oJ;���Ż]l�n>Ai�M�#^��g��9�e�y�W��f���e���䅭�^)���)�X��8�#(}���K��mЃQ��C1{m��bh�-��Mڊ0n�8�Ѹ�f����Py�/4]��u�mSW({hN�П��x�``⼀�P�Q��3�mo�abD&���A��V��;��.^�h�π��A� �r{��U@.�1)�/=}����dŐl���\;-m��1_�Bi�*Ε�����x|���7e�Z������r���?�³{`5���^�[��2�"�4gPE*�Q������OP�1���٫*nي�B���ǰk��!N����T��M��v~?�vV]lf6��`��b�>)�ĕ�̇���n���[v2���/@穃�@V�2��.��,U~�x�CV�rg��C�����ag+H(HKk��O�x�1�U�ϒo��p��U������R�ړF��~*�wW�qj�]O��\������9?����n��
3A�ܔ���W �o�9WN�?�e	+���=��-IV!-���m3o�@�nZXՄ�5���i&�D :��U�3�ԃ�F��`H�nR��n��0��.a=��J�֬�zG����׸�7Zdp,cq�	*�&�f#e+����s��1��#"��"RB3�+݄�>���'�>g�~�k�����M��bt���DQ�@�[2;�6'����r�"��_͵jrpH��*��ٞ%k$�1J\:��Ӕ���=��X���K��m����=�ˤ(`I6�̋t暐�YKϛ'*�"S�M��ڹp����3��|�O��]H�]����k�`bw$�Jy��y����0�~�"N!�mq�DPUw�{Rj�Wh� ����A���Л6;8]<64�T�l�ͬ����F��3a!�#�%�]Vq���Qt�L�D!o8X�g4]��#Y�V����d���gQ��V�֓ԤR���I�h�1Z5Gw�@�U{Vg�ʤ������C~d��)?��/܉�cJ�"MNm6f��R�^�;&��� ٳ�̼?1Q����\�q[/JB�iD�qB�,��î8HD	l��\��J���3�����_�1kn��5bb ��g�����@��9J���iN�
pY��wq@��>�y�1�ۡ��!RH�C���12OudV��ux����F��L�@ˠY���� '�ڐ�^�DY���[s��6�ۮ;/O�<�i��/3�E�続q��m���,�X����ٺ>�5R76HB2t��2z��vYbs��_�f"�d�y�^N������2�&�(3�G�o�+/3�#w2MM��n��x(�P�0�7�ɾ~��A�=]Z:��¦�ȸB�1?��{'_�hݍP���d�Va�ߔ��)@��uP]vf�F#�V����P�Y�0��~Qz��}@oV����=�T������#�.e�M"E2��4>L�Z�fa�B�_��ؓ��k�=C�W=�	�>_6\��]�� �0HO�|�H��uU�.jdĦHb�b.>��dA�l������@�Z��(����=�:熐�@��;�<N_�r��2��2��m��L�cJ�����`G�	�@��T�SY+�7����1;lbu�]Z¶���MY��v��+Xh�$'Iye*��ڦ����Q���!�3v�M�ȏ �g�o'���b;��);lk�\�/��;���O�?!��Bī[۬��Q>w*��q���wU����}OB��QN� &J;�s�$v�GI��#��n��D.� �ݙ9n0�$����@_N�O�`$�-(�fP	�#)�I�������"�cͫ��8i�����k��n4���oV�(?k�h�V)7]�@���>�Iq
ny9Y_�W�,�./��Pvc�����
/�+���QC�!������F���ԕ߷[�S`��6]M��@q;��d	>����\�Y��
(sYZ�� Q��QЛ�0k�2��G(�����1�A�V�`OC!.��*� ���2jdǏ_|c�]su�*qW#��P?3?'3�kZ8Ơ��oe�0���C�D���.�������O]�Wꩨ)q2԰�tP8ð1�^�v�������jkA>?�Y
�\�\��ϓ/��
eT���ګ��̔Ë�W	���˙�٩ ʨ���igd�~�,��@�'�'*��x]R�b�{!ɣc`���A�(n@Dm��/��
vyP�{d�E�W�V�g��	A]ƤIY� ��t=�#���޷=���HN���:+�>���x��L�؛�,��g4��>�$��t��>����o���ڑ<�o"]��ȗ�=��.Qt9	�DۣRԝqv���>�e�o!��ZSXen�i�޽�G�dU`��8�E���)�N�ɝ-�᫽��,�`<�٩��򃚢�"?<��*�P���5AQ\�(CV��@�uW�"R�p�q9X�b'�{%?r�5=�1�JD��N�l���bˑ3��,&�i���=�hPS`�7��6��	�� �n��ȶi��L"50����8�ņ�`޴������m��~��XE�Y7U��(\ը�"�qq�q\���QO��}s�Pl�jHfMa��D����S�2���:x�)C��F������ ��~���}Wa� Y�����-Lsǳ��w��h��]��ċZ8���M��<ؙ�JS��=�F��)��L�􉙘ɺ�Tr/9*�(�˘	�v|���2a?�%���AEM^K�e�*�m*�[o��}.����t�؇�UFq*�`�&��:s��q��]Ŵa/i��X�A�Eoy�/Y���=R~|�e��EPڲ`żY�'Z�d�Ѻt��e�|=h���2�����r�(���8���;��n<��@	0o�Ge�vXy�˯&:a�z�'��X5�̣��i�)q�{���X�($���ea�;�UHb1\|�5�I{��|6�]M��Ĳ����/2��9�U�˪��΃�~"a'5e:j �%/�
}��7��yi{��=�JgC'g�#Vj揹*!m�����U��'���4$��S���ǈ���hZM'�ڄ�օW98�H΁c����0La�fw�1%a�z�v ɞ��þ��qؼ�J
=��m�����P��n.5r��{�����5����RX�=�ax�.�.�!mC� -)1��OH�FVfwP������/���v�TYo]���;�EŇ���fj!,���'���2zp��c�!`�N������]�LǺ��ʆ�G���9���1K���r�.(�v1�>�չ?JI��BRP��\X�ƅ�g;��[�@����	K��K���Iv~���S9�<(\0�K_9��ʹ���
��u؍k/��������Sk�}(v��mCS�ܠ��8-XX|1���R����0��خ��h�	>�f��*��u�lʌx�������V�<��-�ö�a)��<_{C������w&�M@6�`�B�9>x{MG��㺔X9���Wl&	��ք�����U����Z jbXp��.��WA��1u�9��f�0���
S�ݮ�����OS�r��&c��&�d`���Zz�(!�I6dXW����v�k��F"P`��� ����'��zt�(�Or��`�,�'��H�)v)h�~*�KF������c��B�~�Zp�bvV�/��ں�fG�+)�=��#wɇ�h麽��&}�K�;-��WÙ�B6�16Hbt�r����E*��@���tKC'^��4N���c���?"+8	���9lpu����_�L��B��v_Ƚ'i�p���-;X���1%;W���.f@0��8>�����aBE�R���@'t�Di\�p�'����Y���#/%ρ�F�"�+���5:����D�ŀ�6Y�,gW8�;�ĉ�8;T�6���/D��T�]D�,��o����(����!a]���_x��XS����â#OQ� �go���(kr(0g!���-�ĵ>�M�W�AȻd`*�DVK՞�v
.'f(�>yS�xE�_���v��aD_�!��`�N�m��EWb�0��8=���]7���<ηWS��"c��9�fcf[\q�`wg���ZOH)�_�K���·�&M�D��U��XAP���2<y������y$h��"�Zɥk2� �ϗg��_�g�H�u���5�J?M&C9@j8Q�\�Πȴ��kV�"�P���g�z�Uۡ��k��?�
�M�`�b��n����4������L���c��MdI�*�̃-�wǪ�3��C,>B����Yw��G���*f�Lߑ [���V�����W+/��1�J��oq��UST����W3����b �!��M:f鄶~�᫊f�J���?�]�}ܻ��=�^���� 2];T�<dX:QyÑB>*a�hn#��;E)���&fZ�"ޛKX�$�|'9*=fm�L�p�W���˄�a9�h�G���h���+?�c���O�MT�� ǩ��>�6		�����c�nzk�N��#�E��9G58e�~o떄�Ρ�T�KClkMЧ⹻Q���7�6��?�ӑ�j�>)�"P�X�5�����~i����*XLH/�Gӛ�DG��AJg2��k��/����@��I���9�3\�e�`$��H��s��ݦ�����}F��<��v�p��Y�W��ϝ�º�����'� �s�>���c����M�|�69Ӣ��L�Ǔ�O�o9|��Y=as�bY�g��� �O�L��i�U�@���\G�2�h<?f�g�#bLR]:��\�.S��K�9�y�;l'������WJ����3� HO����u-f�� ���,&\ ��z���^UR�$��Kޥn�J���[ڽԎ��l��}�i?�hp�;{-�)���6�Y��B�nZ��@���>��JU�M�
�B�v7��fp�2��O`���uG�G$�X��i�%oT˕��7wt��L���5ء�Dp\��6����>����oJ'a��F�t=P�B�%���|�M=�v�LH�M��R�>���_��L�F�9�΍l1{]Z��V����=/T6�^\�̿n�o������V¦����2�#���*�q,[Ƙ�=��
��i*t��b�R�p=g*[��1�~5i韦Ze��lJ ;���H(����׍�At*��	��%4yRT܉�BI�_~8�2,7��:���4�<ǸU�6��ݤy��:ꅙ�uV7':���DۊR��k	~Xy΢��)
�$�@�֞�U;���K]{�xJTR
˝
��˚(��d� ��&`�����xq�E�Ǿ��K��+�0 ����Z5B�ґ�d|=U�nJ�� ���.�I�Y��Q��10g8��֜Jlb�3&9QLl:8�^-���ϱYxCv�?�bGwB@9�f��5T�;Ϸ �� �gZ�-?D2���!�n�6ƛ����K�>�D�m���������Bل:��i3���#�����m���Wt��7�ۆ�v���^ii�꟣�����1$4�ڦ%�5�'���?ڣ�/�tg<1d��6h��0=�A\,lȚ�����~���@�6�I���Z�a�������S��!6$��9��74�=���M:�����4�cIeru�¨0��.[��ͼ4���9)��� �_N���ut�7��.����x�mN���:e�����Ci�ޚj"��?��3���cj�_������o<`ا~A��N�|�.��:�~���,�<4�\�Hb�l��?�e��w�3f.��x-? �Ұv�Q_��cq�߭��L�ic �ٜ�.ȏ����|����;C��)T���֢����)�Y���{+C^b���u���]��o�öM>Q�"��|w異P�3O|;y�]�I����[��!�I�v��E.���!F$U��� �-y��z-)�o�q޵K���5q�ˠb��;܆w�[k�>A�{[�	���4��,��@?�M��2h���<�=?�u�E�*	�)P�י���@�1�`F�ɠ�V��!UU�2E"�c������Yh�s*�gN��C9�7�a��'>�*W��*��<�Y��r�y"��?׿U�#�s���9b�qFUdV|`�a�h����R��lǕ/\�lǸ=�wr�@�C�8���\��
�s�	
i��F����s���4-�m�.�7H6w~t	��)2~n�Aњs�ۮ�>$����U��%:{gU��G�V�i���w<�j��֏����Ƽy=z���3b��.7ʈ/��aq	+�Hs���l1p����/]��� ]���j����훰Dh�~(���0�5�$A"����4xc���]�H,o�.wR����%_ↁ2߭����M���s�R��\(���eǎ����=��]	��`��
�~�7�$o�0��m��}�Q7e�<�?m�m��
�R��H�&
Q�D^�@?�@ko�̮�O�! D�<�aZ���ƪ��~j�j�`����rS×�T�S���+�4m7���IJ�u{M���9bY���{�{<ڸ��Z��[�P�9=U�̹z
�	�����5�x�v��_ ��_!��,�&& ���P3�%|+uk�	HUyܛ$C��^��yB�ͻ��������8�0�1$�ЪX �bpQ�SnH�d��u+��!a����T��%�C�5c������=��j�i瘿V� :���D_�f����`x��6'S����!}>K/4 b�{E��C~��7�NG)�=���k �o=�G�"C-��;�-�g&����	g�L��Yw&5?��Yx�	/]�P�T�$��-�F0�����|`�"����?�6Z���̯f�![ek�9��V/���x"��T�.{�ﴒ�ay�`���4��V4����핁�߰��^>)�0��i���� �;�q3�D�wi}�~?�.O?�+��me|�}��?D�䪗e@�`K-�9�Wᰜ�h~_d�����pC?{�����C��(�Q�J;�~g\��>j�+��ncj�P��<���j�����xօ�Am���-5d���8�/F@itz^��ar�L�imq�$x��{;�C~l��튋i�v��I�@P��7�W�)����d!������$��S8� �,�># 9,������Ap��cRm��T1�.�:��|;���q]p�@�dyͪE�a����1�N녫��IP���C	��|dPd��;;�9xn$�զ��M�Z�Rc�}���'>�غ��<m��`%79���jq�ű)�'�Ⱔ��7�ayM��̈́�!��Q��%rt�-\�_�hC0���V��8�9)�_���2�[D�e
8g!����'i_aDE�x�)�C<n����A|�*�����G���`\,�8����,��"=�ث����b�yG�@���~��i}sZl;5f�JKI�"�.��M]r��d���c��$�iZy�Qm*���1
SY���5��*OP���	nm���lQRp*R����@^2QAWv�Eg^%���k��n0JE愩��k��K�v�	#��W� u���u���z�;�#��']���)���ΕҨ�8[+�1�#P.�/c8��Zg����������~SZq�&�?��E_��hF,�.��K�ҚP�S��_�}������f��a�w����1ҡR��j���{��Kpv �3�u�OOm��.����]C)��<�.�N<�Мs�>�����֣d
���Dv��u��$�Q�r�.?�����)�y�Z|qLb��o�O����9$l͓_2�7L�}�67���O�����+ƃBH%�y%��jOw��>dpu~�|(�Ά��JxɎ}��kT�)Ԛ�]dƶǸ_KU��w�L����P�-D���(�Pލ� 0G���L�99���G7�}��"���w�3��|W�r�˧
���шD�L�lk�Q��N�(J�jG�ˢ�u泹�[?KH�G�)2�c�N"1O��`$a�oU\�&��U�҇yc�e�*gi��U�����؝>�l4]�� �YX���	����B*e	���_�� �8QV�6D����1T�&��c�h���q�ڂ�1�[i2Z�º��U�%��̈��7ɉ&#N~�]x�o��" �3�������r���B��%��:d�v�������uY�̤����,���_�����г�!�7��� �h��=�G_;=�$b�M��i�����0�d7���?h�Z9
��h[6��HGi{�q`�Wmt�v�<������pӍ p�3wo�7m�[�ގ%q��^��U�FX�A2&�&C��g��ْGg�E�C�qKD��O)��vd��ƨ2����Vt�O��Jj%@V��1	��.�`(��؀^�/�o�M/l�;K��Z �!N�@�8���e'Ŏd/v�}�40�
�t����?f�@wL|�|��=�Գ!��?Z�̹�E�H|\S&�^_Fy�E\�T�d��V3�.;�T��Yν�Ԫ��	�2���Q⏻s��$}9��q:����Vo?m�_J[�܅���%rÉ�@��5tW�0Ա�d�*��"�ut�O
�v�<�Y0Icm�T�a�{���ߣȀ%�5rV	S�5H̉�J!)��p́�t_�e�+wrc��wnѩ���'�)]�2HW���ׅ���i�|��:To� �}��ߜ�0Nz�G��p�f��d},{{��씦S�,�L���ZZ�rb���E��6�����Y���Oa�pVH���vb4bԞ�`X��ub-��c��}hV��	8��������tS9�������z��#�H
��ȕQ��lu6�#�|�%��V3
�R!i�����d,�\�ͻthW� �
z��(Z"�m@!G�&���|@$}��aXT�h�CJe\��dP��:ͭ0A�ž��;�M�E�JX�g�oqx.R�v6����}������\�TE'��4��-�(��3|wo���.>��yE�m��<۟��Ξי}��iX>�痏��?0#������� <<I~�����U�cR�<G�&���)�ʖ6^�T�V���)`���D�`�Q�ȜFX�si�����*Fo 6�@�Yp�È�\=�2⮣)<��ܐ�j��a5�ǿt̚"�μ��%oq�Yx+C���X��B�+��9~���~��`�#�_���,� �Q�N\�\�-��)��3j�v���{���O�dz�&����� �{��_<��P��:��H�s�:��1N��3p���K��$�tU��O6���o�V�3+�t3gH��l��H�����~$ kN܋�߾��CF��5���8��6�վu(#-[��65�Tk���(]�N"_,j2�FBj+a���ܔ3��3䎲,��*�E4�����8<�&m]W��B���R�gT������z��I�ÂڽEVA��5�T�Z�ٍ#�����3�C�ޏՀ�`�J���Z�*��wb��n;�h�ԻR�6g�j{]�E����'�Qu�(���Z2܄qR����눦� k�Z5���Z[l W�Γԝ��P�$4�=�u!��:�N.[iRO^RX�PX��/��-O3}�e����cr��eUv�W+��Ο�RcU�(�i�\W[��`�=J*��b��ؿ�R���Qy:m�B���˦����-I��D�5�LY�:��$�sI��#K���T_�\J��m����&��^h�¨�w% �aص�0��_��aja���؈�8z����"|r)'��ܹK�Gz�
�*C�g0I$�f�YU��Շ^���B����C�t3wmi���ݻ���4����\$�<�^a9*�UF��(�1�>�����J&������x�gg��p_�N����ì������
$��],_3���0���%�3��y�������[�e�2��M�i.*
�C��8�
.�z�����䵓/�(�9�HL��j1�`�c�ʢ��6ϟ��=9Z2U� ܷ��t���K��8+Va1R@�wz�y�~w�8���'7�$�(\]�2��Ŗ!M�P��2^t���oE�}%�PS�[��&rQ���dR��b�ڐ�ֺ0X��KLRG/��z$���:�rd"�b4ܕZ����	��)��� �Y�w.
i��w�J�G�gm1OՃ��N�rK���&�fD�S]e@E�8��-�[g(٧z�r��`�ŗ$�9�Dg���D��|���g{n\��d�|Bhޢ�L{�>ޟUEb���0�-}2vbS?S�L�a�$�����V�򻕲�&]��%��S�@��x��;U��H��콜�����yc���c�� �As<�����nZ!c /�4��S�(��#�S����a���PYz����ʞ�~ʑ�J�|�6��(�{%T��R��`�*{��σ�'lO�V��Y���ed+��9��,�k=}���M�\4�GK��˶<r|mP2n��Ҍ���;�}[�8�E=�(_�q��j�b$q�<}��~�ճ��|�����e�3�r�	N�?��N��s���@�8�M[�=�O�Ds�u��p3��ưk��'��+%f	䭬�7���`���N�����U��;n���k���Q(H���o�,�"Ց��mY�E��
1=�P*s�����_�ף�?�U��m����}�E�6��q�W 5/<Ō�·~�Ϗ��"g�8�������H� ����9��� ���m!?����$|;�$�yο_��0sǌF˷���Ϫ�Z��J�*��6bMιQ[Ӝ����E�}���`�e�	O�HK0Q�
fp���We1Y��� Z9��S8�J��-&�)��cz,����v�!�4�z)��B/�LRų�"�+{�y�q�N��|���$���9��9��rO��i�,{��lE���D��eJ�/-yx�'�%KI��-?Yc���mҕ@�
�0�;��
����:_uJG�r":M�b�o��"����ϼ�� �H2�,�x�U-��IaC�A��Dg��]: N�83ݣ\�p?ݟ(���wg5��`5�i/��͒��Q'�҇�6�F�d/h?�VPpf�%p�)���N˾ �!��f��ʤ{l�����M��-���6�I;d�pR�$bO�b�)�xX*�_�Y�CXǾ�_ɴҽ��d���1U��ε�jY*��k��9��L
Â�3����E�����E�8�Yel���$�XO��eh�v�$7Ma�;�Y-�~�O1v��]L!�W�=C%#P�'>P������֘��H�TqkW=�5rK�<S\��
����˝�o%e��M'�>�G��O�v6��Ƨ>Nd��$D����w�W-�+�E{G�PN̢}"���y�Tu��)M�_��n/r֛gί�������M�U�
�2�c��~*F�]�3��٘�'������e�j��4��e9����fOFB�[>p_���k��͕�!e���A6��t�:�Mݘ�p	<E-K]M^p�!��fp�9��fɞU<F҅�j�M���Wڈ�'�6 '>�Ӕ�T���Q*a�j\h�� mP���e�wA��"�=x�����Z'Ȫ��YJ5>+�`��3B''4�g�
m �S�"�t�o��Ir'�kRF�Nؤ�f��	Aέ<�"� Zcv<Z��W�������)�˸!�֣�>`��z�Ϸ�ɟ��l?��$��������X��!�8���k!��g҇R˝�x,����sOI���E�%�\��G��V���m8Ö��zͼ������6�:2O	M�Xk�
�W�ʸ��l�b ��H��[.��@BȖ���U���
+
�_�˰{	-���6˝��\<C1��+)�_�����$�t[��h��x��੓�2E_�{պo��m�9�X i��c�KAu�:����q(���G�����M��sV����ftO��h��\��tE}!�����"Q�7� �7<W���^�ˁ@��g\����*����C��dD��6���ӯ5�<��4^7^eL���|*�%w���͛LͲ���i?�c!��X�:��t�`,���pi�;����V&���jK�Ē�6Ѽ5�c�> � %1?�������;�O�p�쯼;h/lFz��\F�����Z@fD��DN'NaMڊ���x��L�j�/f��?V��u��������TuR���b	,(9��hB�T�v�̽��5�r_H�@m~�� ��&�*�e��W�7)|�K�\:���(���k�k�+��J�s9a�{/	�M��C�ڃ#�g��1I�G�����t�"$.'��"��,�(����9��>�g����1��OB6dc˖򮿧ܕ\�W ?x)�w	��EP<$i+t�̗�X�H��Cn��r�����}_gH�-�4��k'�L�Mξ�#6�����5`������l�݄�(k-$���G���ҵ9�$��Zb�K��#�p���[�ޕtŶ�/�D�� {5��0U�Tjݗ�����߾=dC��T6r�g�z�}yH��F;d� �8��x�(بX�j=<���2�<}�>���D�3��i�CV�����7'�y�n���#�5� Ur4H��	�L^="`X+a������(��Ѕ4C`j�(5Tb�v�~�gG���Y�?�Mo��j�Nqt��m�6&SVS�ty�8��I�Sv�T�g���P���Y��%�~� ��
���8@���p�g�)�Y/6<ӿg�-{��{��f�HЄ���F�S���X^��QQz�{kc��b��@w��<����n�#;�@�@l{���d�U.\ϩ"T���rH@Tu�je	�2�l����kI�騭�Z|�i���q%бF`��ރʶ�j�M�	)<&o���\��0�eŃo��`m��r�!W! ̐��$���L�D~�,0}�Z{9�ũK	}�]������:#3E=U�4*K� ���_��ު7c�����>��yF�c�D0]rL��ީ��7�����}��5˫�����P���><g)�dz$#2�/�B�lQw`�N�^IK�q�K
��f?��h܅a���{�<��r�c����j���kR:&��#�W���e��n�L�SjCݠ��_�Q��c�:�jdF�(�e��e|^PO�[ъ=�_�>N~U�������~�i������=��!�,4���@(P��|ވ0鲝�I2���~��o�r��c�"1g���M��X�J�eu�g5�/Lͼ>܂���t�{����B���~�������`��̎t-)��p3��L�LB����G�I�'/�rb$��DfQdՋy�\
� �-�0�ĭ�|���^�֖n،�M��~B��k�{�a��U	����5�#�i+T�ʶ�&pYX&X�h�"�O����<�o9k\p������U>�fx6���_d�����/���R!�QL����(�X��mv�E�����va4y�k�*�Ln8�T�(�
�������f/2����@��?�=�fxGj�TU{E�jy�~hD��" ���ܸ\��H�n"�j��&ҳ�S�%)���Ɣؐዘ�m�z��q�7��8����}%g�ICk���"w+L>lo_�1i�������5Fi���ŦЪZ��@�Zڧ5�'ѯ�G�tU�ʺ�V�� �"�gT��w�]دm_��r��@�����ڭ�r��r��V}b���<�jh��bKп߰������"�˿��'����4A9NX�o��z<�v`M=3	뭀A>�,��D���b'��63zf1�W9j�ql�Z��g�`ܻ�i���zh6d52�Ry�F�8�+���3o���������*�J��M
1���t%��~��iʂ�r���N��k��~���
��lĐ��԰�TS�\��h��²��G`��)Y�ٍ�#;��N�Q�a�Z����@d�Y�rb*�~��Gd�hT�u��;v���y(�}F8	�b�`섁�����!B��43̵�1������!��E'�Hk3~d/���cՇ0�#*E��ʃ�!ɗc�9���8$�����iQ?�*ڕ���6]��Ӟ�sv��*��/�N�r�^򑻗&�4�R�&y*���C�8*��u��?M����	�_�Ӎ�(7��p��Ź��t=����C?��%�^@����@�u'م�(-�<������4�ZE��C��Urw�o����|$��H8�<{���T�q6�&�whzy���jEp�՝��	>l�NSj6�nC�5��I��NEh�� �ԬB���a`���k�]j�LV�Q�(n��l�=�q�.�k/��S��U��H������ˑ��/���+T�����0k��,|�tr�W��a�� �WDV �L��)�v��Z���G���A�BY%�Sy���X&�*�?��4�+��S������׽�ŏ�᪦4�c(��D���-S+���ώ�Q�;��N,�4�6E��{Jb5D@�w��^��ѡǠ�MÛ{=ڡ��S/��k�#��3�YW8�K�	ظ��E0�0����jv1���LAP��c��ǿup(�!J [h�TJ�tV#У"8�م]=JkL2�G�G`�U�آ+C�漄�Ė�<��d��=��nk�Fd�R�Z��w���TQ��K;	�}ϱh<�g�&M}�D�_s��p��n�5'�ԏ�۪ H�/��y�K��2U�&~@�����s��!d��!�����P��&e&�r�V��H�M�H~�ZZ������;���ol�p��������s�E�+mbSר��i�Ć��X�߀ے=߶�����B�������^9��G@]bfȉF��#b����v*�烪P}�A����R���	�i�E)1��u��a{�}��g5k{@%.��Pwi�	 �c�\�y֫��m���_Ch��ؿ�Z�X���mLd�SH�B�U??P�R,�؂�j(o(R������N��1e���P��`e����;M-��^���YL�ȡ�&�A�=���}­�;��8�Ц��F�2| �����Z+��L@a��o�:���^IE��A�����е��1�����Q�K��[F����Y@A�i����I+��3f�	��cB����,�]���N8xmǚ��w�~�0J���H�g�Fů�Y�=�9�M���`�X��%����qU�m�,�MH�-��<w	��	c��~K����h/��j9�z����Y{�C���y��I��ɨ������t�j <J@��aj�y�&?��R$X����zq�E��!��p}���.`Z)��6ӏ�ȟM}�T^���F�5���_���G�������6�~�"�D� af�E8� �o+�r %r��� \���a�%��!Z�d�Я���� Q5,�(�+��%"����0,"62�y4�&�f����~P8�ZQS(�h�`�J�q��-��d}�Aw'	΀�����X�v�
Dc&�31���[Ҡq	kjF���1����K�,�O�����X�X�J\��hF������W�V6�գ
N���:o���a	jT�L��������,}�QKj�'W7R�!z��9mK\�	AbT>�r����O���7��k��1R3Gj���mϢ�O��
�0�+t�3h�;�h�Е���~8��z�@U:Q���)��ya��*�v��h���}"j�"Vi|o�/4�=����a=D�Mֵ��G;r�T�?���e%�M�Aq��	
��K���L��ɮ.\]��;��
Etv�QM(����^��ϋ�j��[*1��ت�;�x�W���p�@S*%���"I��*�4n��pM�(e�ݱ�U����c+����(~��d���+��#S�3�ވC�]|�����$0H�$�盐r'0�����R�!�~v�|*7�a��N��pr��&���T�i�e��k��Ts��&���z:��@��F�O.���M��2\�Ρ�B
�|-'�'�e+��
hO7��L�]����f���D|����W�I\�jܨ��� �k�H�j��Q�c��f�y�XEҲx\BHT{]\�H�R�M ���G��Oz�z���.|`��b|��,w$@**�1݋��N��N��9��P�+���_2R`��ś�mȥ��3�wWZ������F�{w�@dhbg|��	���a��Ԣ<���G��[�' ��S~��c�M7֯�ԁ+����;�mR>���.���*�/�&�w.=Z��i���cKY賍䛒�������ӷ�_H����L�KI��<B����D*�d3�G@k�n�=����~���wa%������OQ_/�/��J/�}��V$�TK���K��˷�9�B�
�vF�m��� nް!Ա@��N*�"ƠJ��F�0K��b��F�ٜӨ%-��H��߫m�qLJ��ɖ��lq��7<������(�(}tu�:�}��hLHϫo5���z&�������B��(xY��Jd�����jU�d���z��/�-A�1�݄���s��7Y>���]T��[#/w����v��i�,Du*�M_�k�i�蒕M~��(nSR������Ǔ2���d�-&F5R��?�5=�6D��ﺊUh?��<�B�}Š-&z�[߳�+�}�����#N��N�X���ґ`c�X�zR�Ժ�+no��Ou�]mGu��7B����6b����^�q���(N<�������ڿ�9���/F8nQz	4~e]Xhě� ;@��4N˒R�}�ͨܔ+�� '�26k]P)��ζ��{�����X{_Ҫ�짎MF"��4R���b��~�ӊL����(���/�Q��u�p7r��7���;���q�b�rֱ�2�t��c��"������F �G�4���)V�v�"\�shWҁv6	��_/��)#{���ĥo�X�o�e_OvMo,�:΅�J�l˱��"�N[��a'"<�;"vR)��'5L����f��rgG �_ �T�	m|�밫 x>�1oSOKh��{x���d�2�|��Dc�b�B|��\&Vx%�dr9��K��^���3G�r�0t�U��FF�>�6F�Z�0��3 �3����]3q�
�+�+;�S
o�Ӟ�5.v�.b�:�jl/��V���a�\y1��a2S��_�����(^�_tQ�K�J�5�s�#�M��<����|k��F*i�j�3�<��"���1��8_E6<Q��Z9x�!0k?��#'&�v�;P��-�Dr2�9�!���/�N$��\� d^��m)N���Ḓi�u�ؘ�%rߪ:"��H���ub��*��2~ȣ�i�uƎ��&�l���+#⩪��H��O*�������VZ�	���>�j�eib�C�4�҉}�85�q�ߣR�\?bp�%Jk*�q)�B�CP��|�ptw�6��[����U;������9����Z%��P�fi����4+�;�@�����{f��^k��_�%���	����c�Q	�T�
�g2����ځ��ƿc���87�����\K�>�1z��*��`ў��[vT�Q�:�hd�`he����n�[�%ܵ�l��ن}eY1�ٍ ���m�+����Q��H��F
4p��7g�K���fT��94֭�;����)j���&����������Y�V|���B�y堢�}�q��(���O�As�}C�7�J�a_��F��[I�we��^�-c���=����1k�B�v�֔��kL��W��iO�r��yA�6zn�8%Z�@W��a��ف$`�7�R����´D�M>�vƂO���UʔH�����ԋ[|#H`��f�3��
�7���;�D��FM�!�~��2�R�D>���^u����3�K*J���,D��5�%$9G��$�7l��wy�� �y���9�o�W��I����v�*T���qv^�����L߅V����N�Q��.{����)�:8���{!؃&6�vZ4B9����E<ډ	D_���NdO�i�F�}Ж��FJ�	����������|�q@or�H�
�%��hds.o�vL&���2(�T��xf��2Y�d�h�t�5��Ty�����v�I�P��)\6pV�nx� ^�.���BZ�U%��y$��CQË�>4J2���kXlܘ3��a��$�s�������z�Ƈ�爡�Xx	^��d݅+�P��M�Q��Ν�mřx倍8�Ln���G��C�ءa����c�S*"6���㳑���$7��a��>^��6�a�.%�����Bc���gn$j�!�����ƹM>:���;�\�*$�F����EI����צ��Pe��<�V:A��>�U��}3m������p��036w���7�)��#��U��LQ� LY8��yZ$��Y�SÑ4�Ό6$��:Hh��Ը�!���}_~Ls�� ���s��3*&YD$�ͻݦ�TP��jM�͏�Ý/��ߓS_�ɏ`�����Cs�k�8IaKΫ�|�u�<�}�KJDS@�e|u?/�	��Q�����#�P���I?��O����!!7���Gd�qH�O����������yʺ��`�h����>X�խL��+YO#v�v���:�vp����*MVB�?"T������gp��r�'��Q�j��`�kn��^v��/��3(�#���n�#����m-b _C�����"��6����~����l�X��h|�@�xҏ���׋��é=��
-�$Nx��qq��V����PzJK��Z�#����vW-:�^�6X�W���(t���+�F6@����g�.��tC,�	���K���Eî�;A��Zf�n��= Ps�-�\���?ŧ�֖�{Ġ
�y�A�f��W�4�ӳz5�z�:LH�_�o��CG�9sKI4��Rǒ��
�_z��]w����W���ǲ#ԯ���x���p�<$��67���ґKJ��Tw~�Nl�՞�F���h�6/��# iƋ��o���E�p�5�h􍏺���O��փ��J=�o����ߢ���c�"��
,�΢�<A�P#�?�K�©������O�kg?����y.q�D@?�Ǡa6K|,�5�`��/
�U���(B�@�`z�Z��q��oX�G]�-YO�ici5T���,�FA�MV6��i6f}V�M)W��;�_��#��GK#��_E�Ж����l��v�C��K,���h��0��[��SVhס�0��`Mk� .Ը��θ�a����?vx��4}@�uS���D�7̎h83�>�_9d���2�!Ʉr'G�ַ��K��Y�[�dp�*�>+�ty������Mh����0�p�A��a��d{"�P����[� ��>-���N��U,����W�1��ڔ�6d����=�%�� ]A��|�����4e�3�=d��9��"xr��&�M���kF4����C��8����~!�Ҽ+5��(�%��W���޴?&sk���6��=��(�u�����Tq���vwW��$2�d��5��jw
���\]��yo��1)*u��iqt�b�.�b�)��B摻���ƣq.�{v�9�/�c!!�l?F7���P[����J��k,�g䠑�w�**tӅ����5�k_7��Ε�Q��o����,-� �d;���1�0T�T�]d�mk���Y��D:h�N���݊F�F:o�V�}�l5�̸�'��G���=�#��J4^sׅ�q�';{J��a��2���r�C�2{Ԑ�'��8Ct��$���p-�򭝻���8x��mP����Хm�U�S��
�^�\��m�����2(�et`_�/8��@�m�=9���Ĳ�Fxsc}��Ѩ��X�j��r�_�|w�S�@��.�"%�izU�s�àgL� ��=����B��(��^b��p���o���,AAS����M����#�<)혇>^�6N�q���j�C��|�[�;��C"A��A��/`����D����w��l�� ~�),�^λ �翌gA>���a;+R�lds'����;@0�c�q�z������Z@��\�]���οI�ٜ<.z@|8�R��H�dG�b�Eҧ��r����%�E�v�P�}f��X�J�K{�~��<���ρ���/4ȎE��N��X�i��N7�Na���8�(`kP�b6x��-��X<߽ lk�~�b�0�-Z��TQ �&�1Vo��kk���t�s����e'`j�y�G&���C	��E��S"P͖���~H߮k�ç#� g�Ϗ��%���|g�K�|��)�,o)��ڃ::Wد���AWL��r����޽7��#M�G����F���~��I�̰��U�|ֺDY:a���r�T�j��k֝w1sħ������\')iE'�oLE������7�.�+���L�	_�x���-��D0��pI�I���E�d���!�c'���/"Bb����Z
��ʌJA�*nrz�)Y�E�:D��݇� �A{���f�n�q�-�c�� �,�C=y1~�i�(�M�&��'�!���b�}���
���ͦnvv��D̙w�ӺCuˮ��b'��+>f�9��V?���>a_����,�ٹu�=��#�|�}3��d�0��Qo��cz`�X��e�
��e����,��ζ�J��b-��8�:�� ��/T�a���e�!$p�!F�<�~U2i\y�;l�)j�߶
���*�Y񎃅��ʍ��*�h�X��jU#�WX�B0�����U���a>����.�E?�ڽX�R��_uB\��`����9�g�kFU@�<2E<}�㕮�iє��5	o,W�,eQ�~�}ƛ|E�w���k�+�#����rt4�1�-p�m۽ٶI~��qx�`9�bG S�W4xr0R���M0F�&čtf�f��3�hG����EsC����Wy��Q$�q@�xP�)�O/،� ��ha��9q�g2�^Ұ���l��J���$�щ��3����v��'�d��[5����ʅ�f+tK2���"'����?�!7Ġ~�y��q���_���Ohn}��&�%�'���C�{�?9e���� ����ѭ�D-8��gW��� B��M��1���n�w������9�ܝޫ��h���3V���7�<��F>�Z�(�g�g U�
�8ʎ�Q�W���l��վ��_fn�������|,�݇u+@|&�5PU��TQ���I��?���� ��G+�qL-�J�h�疢z��T*Ut�'_��-_ծ����@[�yWƐ�T�֤:te
�,3�MY���M�!�|��Ĕ�ܶ	4�7��u+'�Q��)��&��ݼ�*<l��-5Rk�$�Ѥ�|zw�^e��e�j2RG����F5'qu�u��W=�H����f�=/�6�V��LTh��7�	Y�~��8A΀��Ɋ�4_�f��@���C��:�w/�`g��Պ�AXg����E��0��X,ӿ6�k� �����������iH� ����p 3� `��Ѓ�Qv��}��Z���3[�8R���؅�;=ϝy[ RI����S΋�4f�VN0�=�p�}}����h�on��^qCO���gnW)�*�:��K�r}iI * �&u�(�H,�5��5P]����)D?�Gm)ѝ�A��� d�Z�7���d݃�@���b��̪C�К�Wl��6s;.��q���U��c������ZZjoN��?XȮ�dz��?2�/DǓf���R�%<�j%h�$����S�yȜ�m~��Ga1���V,��n��J�V��`�w�j?7V����/�CN��4ԃ#��ۛgj��n��8s�yn~C/+y�sD��k����zm(�x���
o��s}��>�.>;Z
��@QT�>a:��Z�������Ф�N瓙�Y�c�9_��Sʝ�9.6�X�_V=q�B7xC*�i���
L-Ch/j�Y#G#����D��]��8�-��L��6����|6�>y����uE+O�B{�$�����vZ"��̗;�nf��:��Hz�B3W	�9CZ+��I�u�u���&ӏA���3��)QN�L����?IJMH�UHsI �Fl!�u��#3��vwP����-�r�[�I������Ò��_w�Ain\�+��|�E���ؑ��5�l4u�S�5s�IQ�}O���9���	��v'��(G7R��҂%��H�-U(�I2�=Q�	: @E�����Y(6�)MF��5��Y)����]_�d���@��?2�撩t�&�%�6*����q�����H{<I��Wq����ʴ�9wEba}q���' '3 �̶��� ��3}��J�Ƚ<Ю�.�ػ���+(,�hi�S�d0��A� cT��`K��tF*�s���I����V�y3�l�Ip2�E�����`�m��pL��������V�?����
�:��,�f�X�Bhw�pv�ڤT�P�p��>��ھ�sr���c���
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�쑃)�˴�V����u~�@���eUf��8��ַ�l|'|X�
UI/nVK�p�gC�3ʵ�/yz�"|��8n;�e=b�?�[b����do{��%�e0������,�CDS�H?�΄c"��M����f5�c���Ц��G�i��~ e�iE��;��s��}�|�;wa��Lh����-��J��K֜(7G��/R�1�*����?�=����&�]:,K2��܄h)�^�+5��?׵n��׺^N=�jL�\�W;#�qT��+���%��,Ծ �S���A�C�5����]�x9P|�r�;���h�?{�D��v!4��x�>�?5���k��>8��y\.����W��]�ͷ
V�i\zb6�8.C���X)d�\����xj$��MD������wZ�򐸬FXP����M��`t����U:яP�exj�)�_M{�1p2����s��5�Nv
��2�8?oD%��Nӑ�u�#IEd����hT���q���`	��F:]�u�}��L�>�9������Z��^�
�.�K���� Fս��i<;����Z��\nZmWYd?�)�0�f��HU2�7�*M5T���癦㸶ZcD���w(�����'�&Á<G��6�	��>��7?�^�}C6�})9�/�o�Nv�~�<x^�[�d�I�Cm}���(�ݺZ���8�~K�W�w!8�QT/�wՈt�&�Âo�K�v��C��H��U�|�Տ�j�o��j��4����[�a�]c������q��k����E�΍�Xh�.w��p�B���6n��S�6:T��k&�7����,g������I��������:9f���U��}R�`]�ZE��I�]7���O
M�Z���O�zl�L�q!S�ث�O�%�NJ \�aT��r����c��-,̶ۖN� gRt����'�%%�FT�k�o6� S,�[W%�n�r�p�����ݵ��y�".���>Zg�2m7a.`���d̃f�
\��{�Z_�xǟﶊe���YL��l�q�s^��A*g�LT�	��d�C�P���[ɸh���~�b"N��D�Y��^}�t%����i�=�G�P�!t�ƕY$5;$�9q<�_�Ӥ��Ĉ�Z��� �рb���q�X��;���#N�F
��*7�9�z��<�藟J㪃Ν�u=$�~g�D�"�$bjc�����Xs�>K��G��[	?�Ųͨ�jp���:�X���T+��r��O�4I�g�S���v�	Y<�wY��U�)+�<F)�F�����������ʫ��b�*�
�F�;֫Eŉ���Ho�HFH����b[��p�r��;���Ui۷i;tÑ #�slC�����Kq߃���.�v]K�pvx���8Cx�q<0���L�N�G����ڊާ��]qkv>I�)!�������[ �G���A�@3=r&z9�]hk��gr��6r����@J��D7/��0a���VZ�<�@Z�z�%�ިND%|}ȌV�_ڕE��������W2!zq���՝�ģ=V���}�|��7J�;�~p�Y�G�*p�b6�o}!s��b�5�&��6��DV��>��4-�����
W � {�G��ƌ$"]���U���=���ߵ�!J���8^���a��p�+�[+����龎K���u�3egi���)P��ի��it����o�uu�����\iLk<nK\5�zU�F�w���e�	��p�3��^��M�hI��<�:fpݗ?�~��b�*�f���@�<�A�V�f`!z�&�l��2��H<BV�z�m� �/��X���9�'��4�g���S�մ�����B�.f�7�W��"�6f�LmpK:AX"�y��`.�~�	\)C���G�/p�
_�n6��ˏU�M��B�>�HW ������Y��w*�3�?^�x|p�0�L^P�_� ��	駦�=�ޝS��h���;��呿ہ`j��>"�'�xQA�M2��l^�E<&��w1�l
`��3^������)GA�V���k��\�Q���Q��NLe�3s},�3Rc�]T��j��c�f���e���!�yQ=
�� K��)���t�O���n����"Ք�
�M�<�Y��X�����Ƥ(�S_��Tb��Z�vk#ߢV��6*���v�BY��q=J��*��j5M�-WE&�;�z�"�b�D��T����E�G,�����������`HJ
N��X��ޞ��X��Օ�����am�M�"k~;)��+)>yk�m��%H>�!W:�No�F�����A��<Y̆�mA��U�|����t+�hLO�B!���&�D�w��jI$i�$���K^C�c��hS��"࿻�1�Ck�Q��5M	sX�v`��.��'.d0���?���2��C��O|��I�kb���(��O]��G��)�4�`?�F!��^f��G���Xss�_����AR�A��<$�����D���$���� �V�=�T(��9�R�D���C�,��� vy�ߵ�쫱�ظ+���4��c�Ϊ<�|�1q�OEmg�:5�6I��6`�	l~%�<�@���v�b}��a���7S�w>��i�U``1����H�����q2v%�@/(8�[u`pHX�2@���F�.���Y����|4(�^u�>������f��c��\6���(=N��/BD�#E5�a�>�Κ�<� ݼ�Q���\8�ͣ?SH�3�vFRX ��]���O��=�	��k����,���6�YQ�0�n ����g��19��"��fwpW�����q � fS�7���9ߗ=��WXmc�>PH�+�%��J������Kу���z	2�~�{#$ I��%����p��r[~ō3uøM ��|�d�Q:}J+{���w���g���_o���Mp�<>��O�����_�0�9���)u�_��?��݀r��^J�L&>��I���6o0K�S���e:8�{ASp��#������ @�􇦍O��k����}D��;tlYa("�Wc{ �b=��in���<�Z�e>Hi�|�F+��P��>4G�x�t0{��w���'�+�DDO~��J'nʈ�"��rU��:Do��Ta���&��-t>�t���[0�|XG=ݭ����V�|l�H���z�����B��8v���M��4n���^��rrk�����<Nx�q|������t��֐��'�Din�Y�|��#,��e,�q쥍tQ����W�;"�V�ʩ�e��~�����NCª�F5�<HVck��9���_	�5��~k�"E<�V�"��%�o��B�IR�HKћe	I�4����j��u���fa���lH�G+�A�����H����aR���P� *sO��O���r�q�͚��f����z�4ݰf����Do��bWDf[�$��{ec�S��C��a;����۳�V=���)�S�+�tuXpX�oH������S��I��<5-˱�,���V
A������*��r�d)Mz��p}ӳe_e�k�eXA�>�v��b���q�5�|g��mM};�R�Ϣ F��s"�C�[�\C�VQ��Ҷ���K�ҙ�!q.**���)NV�}(G����X/�aQ� �1���O�/_��H ,�L��/��L���ׅR-��:+*��ʭ�fΠ_������H̅�ɠ���x�*�u�un�xl��ȹ�����z�ÀuS��ʷ�W������x��c���1�_k�@U�he�ȼmRI�;�j��5��XBV'�
A>/iG��p=m-#z\�L���pT��A](�܁��2�h+�Q�Y�;�H���D�`��:���dj���^�|H�H֡?w�4���fW���oc�m�;���]q!�8{�X(�C
�$?�����j�^�oP3���7�SL��S/w�>���V~�AN����ȁ�Y���P��W@<��{_��gĢ�]2�/G1]>��vW[ī�дN}E! �`+2��3b�J�w�
tC���yMǱ�eu�09S)*."@���tI�Vc[g�3���	3j�K������)�T��059��/��\C	������9̱ )���
oi�H́tQMU#7�8]!RT����+qK����v����O�w�k
�����~��A���w�;Nbq}�?�*�����C���:|��O�B@q-ߜ���aBP$o&v�C}c6�^P��kq��n�D�����e��*b�N��c��UdlW4����#��q���������k�a�k̏P�$&�W��2�_a��(L`3Z�@{ߑaC�T��O֟��o����`�T��s|UL��_~٪%L�byKMjK$�m��-I���Ͽ1,1X2��U�
59� �����۽Ue�=�S�a,r�o���F\Z���~��Y��j��iT>���� *�9���t?̖r�P�	o�5����Go� MIE�״m4�8Ȯ*gCpV�گR0�!�	� �
���%B�Ϯ��A���2T.pۼV�`�qȑ�b��]h#�Ϡv�7q���!��.�3�<Սv�/��g��}���5��&2,`F(�/�͗[�w�FvB�q�*-v Q�˨��&�ܯ����&S����#B�k�iU�%�w�;b��4�i]�<���������ƙ<I�;��%��BCr�Cun�4$�3�M^���ް�Ә�>���i�OPBcL�֮�<�N���I,�c�e���E��P�M�'����-���{�y�4���`M�:��_�(P�W�BvBJi��S�&Ks����1���`o�A�126�퍽�wmlV�mH���tt��m�������J1,�@'ȑa�,
���B�U�Z!��=q �Ǘ�P�۫,�ʨ�Ɋ2�:�x��������d�g��S�s>y�)�����Ò�76�{� "�W1��6
$��?d��%TlTD����`Ml�=��62�M�i8��;���NO؅(� /%VU�� ;'.$�P���B����iG���3�n�p_�@h5�rp	ш��}����u�BC�/*Xf��w���A�q%F��H)W�ue{%{��M*�X�@�KM���&�1cl\I�*�P���d~��TA.'�����Aۤ�)Yz��s*�L�a����$�8(cಕ��{�0w@��%��I�g*^�R�ף�̈�W i.�	SG`H�s� ���������.�ͩ"wS(�c?�����y.:���+c�W¼�řɉM��͹'��~�:�Ϲ{=X��?u��ь�
��A��j};G8,�:���>o��H�hA��O����Tdh�~��q��owF*cr�>`�;��5F��y���`���c�FVyH���rW9alSbr���(=�:~��W�v�[���2�C��w|
�.���H����K��9�o��]�^��fU�?�Y���3i�lȼ5��8y�s|�p�����2Y���i��Ra�({vo�ys����)��{�N�%�{���K��V�#;Pr$�,f���O������$��e/��Ağ�X��k<��W٠�0��g��)i �ܮG���db�aϞќ'ȧNJnJ̑��8Fs
�sGG�Ȼ[��+Ը9�f�%,_��{�]k����3Ѝ�j�n��J��$r��=���*Dc�����ŗ'=�����a��D���vH���C='�`N�gt8�ݤ��&�ƒU5�'�&�c��@�y��׻�5B ��wWs��t)t���
	XT-~w��IN��u��C^3�܁<�=(��E�h��Rs.�zT�FTCP�f��Գ����Xp����Ԫ���AK���$<����Ƽ���b��5^Y����쁾���4�/ehy�
��6�p�5,/Ή��6�I�?��>�W�\u��M"O��P薥V{�����^2���޳y^DC�R��Aw���u9��|�5��6K�E�J����yV��kZ�C�m�=�8�S[0�'a�k�.V4���lZ��H����8&IU3�yE�x/����N��Ӡ���dth�8u�䞕�Q�c���U감U`<��LQ02��_P�,uҒ17l{�1�f�V�&p������st�����Y1,r^�T��f��Uc'��)0��*�$m�3��� ]\��3(�y�eZM�4��A5W��Ҕ���
��5�z�ǖD�T6\�.X�Yif�,9��)�6�4���ӑ�����7��N�5,�E��STd`��PF#k�vk	ȺxF�j=���*D�M�#nX0+
zp͹���Af�ek]{����_�� f��S�MGm玲�Wy�Eb~���38�0��	 ����&��@�!��5�i��|7�1Sf8A�]�ޞ��^[���s�磪�iؤi��ELx��sXJ�8��_5Z�Q�-�]G���4��e�2�3��iD�q3��ƀ�XK���OEe�������L�-���>Ϭ��i���uש��Svgj�_�����(8}�gC�OD�}�C�oqݟ��� �P��nF���[��*j�o�v��=(M�fCi�'s��vz'���^HH���ܤ�f�m��/�U:-r�^%*�m�I�6����̞7y�:������8��@ⴛ^�(	I0N�i\<��'���.s���>��Sr�q�H0�h�^�k���9z�f�Eݴ���N��ug�-�Ṷ�vR��Z���&4��	n!���'"��{DO���Q���z��Iư�K�C�r�x��I�jV�_�ťƗ���۴�^l<��%x��m�^/%0���_�3��i����R�1g:�jQT��r���KD��*��t49O��I6��	�L�0�zb�Pvr��.��'b�ț�vrn)��a8>�Q ���t9:�������&y�9D��]���;.S��oFH���+C����2��ܧ�8�/�`�s�zQC.�L,�9��p�ۦ��ʙZ���?��G�:�f�w��Va���4�zwHVooP�$��w3<��
(���|��4�80�����p`'��,�У���#���/c/6������Bg�E��p<�Z�9�x�>A �G�a��et�k��q��(�J��@�N�F�M�`���]��,�����f��Π5��h�����\9���q���-s�>4oC7(�0�Уl�(
�f��X[�4���*�y��~���rZ�Q�{�}��_�[�u��6�J%��&8�������ƞ�����$}���p2sk��e6jSZ����!�"�|�����a�~Q�"��R� @�[� $�<��ڄ�[u#���GK�$�2�6��}��y;C�d�?�v3�K��(�%� U��lx)MD�OE�X���zi_����i� α3�����ʄ���Ί�b_����B��ʛ����i�dy�ãr]7�Y���.T�\�ר� ��@-�r_i�8R��أ#�N�*�v`8U6�_�i�w0u8H��w�����RT��*tZ�w�?6�1K�^Z�^�P�d�Ǻ&���$��q$��o�>��+�1Vͱd���gw�.�0�A����B>Bvv�ʛz����wl�椚����BP�Y=�"n�fx)��%��O�����ӱ�rK*���D��Ll��נ�4c5�9�]��E-ҙ�M��ag�M����r4���<��` ojҥ�~���ȼ\*8h	�_�O���s��� �<Ɲ�^�9���d�WU��qemDW���x�cn��,%%�v��(a�[��;o��\z����m�����B�G:�>;:k-9D��܊�K G`(1gU(/��j���)��,u󒔵�ۮv��n&Úc3�,�kR��Q8̘3fP���i8=����])�2��f���6
�Z�J
��bw�y����,ښBf0��i�����a��$���4h��i�<	�9>J:�dح9K�DgD �~8���u(��{��aZ�ω�}��&��À���z�2d�~z�=�>YE1�wC�w�Q�[f���_u�*�#2c�
jNF	vP|)��0�s�Y�{(&;�#��$&��ewK�����?�ĳ��;F_�aWR�=��n�Y�������4�{Np|Yl_a?Q(�#��>W?���y>HT�֬�.�q�P�V]�y�ސ�b���L�i~{Ď���	a��)ㅩ�4�����b�rK:��TYO���`0�l&M������Ƌ����˾�X�a�>;��S�;����2ڇ�>I2q%��xǤ,�� ¬8�5��{=���w��"-��ma*�#*��z��i���9���o�~�������s�����aL��-�gVݠz.
L��bcelak�ee� 7s�k�턀�"+�T9�~�"/ȹf��b�6���w�u|�#�&�.Ҹ��z�R�&�`)���p�מT����p�-�:Q`��,�L upбl�!�M� �x����(F�J�R-���K-&���� ޣ��+������t ���f���Y>0o�����$�`4�t^x���EhB�Y�����϶��_��a�l�#��)+�T�OJ�	0j�H�!�� ډ�X�O=�#���Gg���A#���.�͝B��"C� ��n�������0A�Q��,LP�1�<�ٮ����3kq��ƑD��w����W���N����ߛ�3�i���|(�� Swj�š`�����7NS��V���m�F1�^��r����NJ�}��c���<�C���- S҂�E�G	�$�A	�nŏ�Kp0YgE9�B�� <�\X?�V�?�h��a0A��@�G}+6���'���$<Z�R���n�߁䷴b�`�vI:�m�����&��"�y
� ���K�w)LP(��2k�}A勼)��A�7Eܮ"<[� n��h�z+XQ��D1�!V��d3#��g�|>���PY��@*�����ɓ��L#ŀQ���Y;J��!�w�.N�A`t׻x�T���51���(��\"Xb�`[L�H�ZWҦ>�%et��՗c��/�of�Xr�?Ӷ�!��Z�ڂ�*�7�(aHj����(�?B� X���ޜvaY/�d)�u%0�!D���$?�e9�G����6��E��?�z���N �bs�)!
�J�~�Fފ�`��CDv;.}��yL_�MY�G<e�I�����jis�`vA���%o8�c@�x0^F>,hmJ|;���Z�;�<�4J8	ڃ�r��y�2��٭-�s3U5U2�(ئ����q���1u��W��rŀ��_K�iCY�$��=Hu꽞ܞ���@U �ɐiӵ9I SO&<LS��X��jq���\�g���4EPbĠ1�sҽ߹0g�E��K�3Y��#��Q����	�S]���U��&��|�{�����t�7[�6�S/-M+E6P�@���0���%���'m.sP%��I��,?�����ײ��2$������ȋ�p�̡+H�Z<<��Es�. �,����rƹ���4Կ-L�RNL^g|�R:� ЮR����7�'DP��Uyx�k?�Q��������#c\�|9qg~ƍyS�5��
}:�<r���aOb�����`�[�;�y[b\�i�#��Q2����[��+�k�T`�H'�g�X�	������+k�U��mY�t�}�إ�₸�%kD9���>@�"&�YTp�&��r�/�[/8�ͲCЗ��T��I�_�b&��-\=��W��b���(���d��D�?+u,�5����gљ�9� ���O��Z�AkY�Q�Z������F��(� }��ϴ%"���퐟,9�E|F�	<G��w�?m�ư�R��ةq\n�[J���8YFw�p����-�XiX(�ES��]��H*b��~Hr�	� ͊�x6���)��Z�Y����R��2&v���D�U��L`)6A�>o�x^E��vl;��й|S�r��sLڋ`ml���p&2x3�:����M4�Sx;a�L��g���w����\`�}�'�Ɠ��69)3�0A�9��0��/���GN��+�q_~�7b�5�օ�e�깳0,3Δ��	�����
�ɔ�b�{���8#vT�Lq�*�����]���8b����d�s�ؿ&��5����J�1�!�fK*i�g���sA��f���L��i����<O�o4��J�e�2�t���#��[�~Z�_�H֟>m�:�Ӄ>�,|�70zT�����'����BI�h�@��U�?N[/ר�ƹT�=��˽?2m#x3 {�=�5U�0�����n�!\E�
[7m
s�+���Ǯ?���ҋ���%INW��A{�d������ٺ; ����`��<�о��i��E5{�R\�lj���f)˅}Ŕ��N+n	�.��$���j>�.��$�'�u��T}"� ��緖B.�Ix�v�E�^a���(��[��t>���M!�<y�\�E��7ē-L��1��B�ղ��n����qK���9��3��1����_�H��Jy-A�d�6��f ��z�}jH,����n�؝$��������=�r�:
�e�Y�򵍮:��
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���|���t�9?T�]'�=Ө��B.8��k�����F^yW#��������3�����W�\��U�mI5�#��A��K���A��]�A����?����:*�+!8j����rb�Mm�6��퟇�1��忥VD�,�*��sgI�%�1?���p�hP���8+DE+4��
*��i���� P[:_s��&O���b�������Fu8iZ��>��U3��G��'�2���nq��K�0��P�ou��UDneNNĒ`�'?2�6���Z��}jEt^jH�c�Po��E�NA?��X�̇9}Vf�]������1FRo�[�ch ��*��_�ҳ8� 0��퇛��Ò��PucLԽ����ԙ؂�{햋i��������5�2H$�,���JTѶ@�Zǲ�f���%��0�ޖ�'��F_�A��uf]Y Pq���3<wO���#x'������*�͎Eoa"�G����K�-�Ϲ��4����H�T:��	-N�Hn�M��GY���I�����T� ���A��+�e1�]E񹼷���M��Y��AU'v�b�l�kb�6�a�!G/AJR�xo1Ur;��N��p����&j�ibp�U�&)gP��[��9���zJY�-3}!��MT�Ev�δo(��e&���E�a���uC�E+�v�c1���g���"�YV�
�]|�.�c河Y��ݤ��Y���c23�����r��(��( ��-*���-������n�5]OC����3L0�G�]}�$�̥Uhb���oG.�:��vWAa�F:��S=�R��aە2<���	��N�^W�^H��t,����y�����2%ir�-)���#ʂ�$�k7;��ֿ�'���۬�v���_�ne���[Tm��jD	���?_l��7��T%���2��=ȝWrS��qY�u{�������?�7"�Ipo�H�����8,K��;�r]"��a����{Wk=H�-�R�+��nVJ�� ׅ�GE�@���TW�ѽgg�E�EދC(�����vx:/��r3��Χ�j��H5~_X� ��f��$��ܙ��gI7����4�:���w//�.�I�:��N����s�π:r�m���5�-䳣I��)Jי�>������H �T8лc�%RƢ��	��q�8������P1xpꕆoؗ6��ST��_s(�v������� ��L{� �sA=_���8�U�<$�*��&u/^!ܔ���yHy�6q�x�ʑ�����&"�5���Q�e���4z>�L#UV!��
�[�����v����O��f�z�_���K�����5�?g�;�˽Z���Ր�|q����U؋� l�r��u�tHX��|Ssy���=C�q0%/+��}#�&,���뒝ʢ�Vw�Q[�e�fq�PYd�*�¼�`e�3{COԢ3Km����%l��]~��I
4؋�X�S�m+�h�ʀ�FTT�F�qx"�K%�!��D*g�ZڤY��`��S�������T��|�[���JN���?��a�p!u?tY��1���*W�;�����(4D�G�":tyU���R#K�lf�J�7��S��|M���z����,�o��P��R�4K)3��_�����2N�Ev�^��_��$���НN3=��m��
�G � 4K��˗�3:|]43
�Yc��U�Û��Ui��=�Ôp�7`;S�g�.�g\�c�	��,#;�g PR.1�l'2�_]��N�<m��y5�>�bA���+�R�.�f�=�����.�h�lSL�m���[i��p��A\�L<A� lc?)Ez~��ڽ�����%8��.h�4A���x���C��M@�f��(���Vn0�� rQ{U�[���)\,�69�&��a�Hp�u��u�,ū�@<9��߻���[�v=O=�����!�OOy�;���"����F����X��U�y��c処O�^�aCJA��`f�s&���K-��Ydp���%�an��1eZl��	prx� rf[?���B�w�#�R�ݳ0?ÜU��p�\d&>�N\(�a���H{B�-/�o*�@�?�kT�qC/>ٝ@�ʍ�/W�Hg�/�F��7�z\�1A@��ut�j�tg,#��r�����tB��%�}sN� ��9u�֗h�J���^^�G�'߄�ܘ!�OŠ�3u52H�]�*��"kY��:��C�9��R��]���:D�>��i�[u�j�-�+cx��BD��+���J!z*��nrnI��Z����}�ñh{���� ��UЄ+rR?���+$X�4\U:7��O�z�䕕�^�����~���m�ba�O�����_'wM^w�ާQUD�J�͗��g$�b!�5Q�L`�cx<�L����) �P���_�>��6r�w�͘D��9��|��愗���r��?�*a�7�(�5��]rk���a9B����N���r<aE�8Ḫ��yt)H�Id	�sn�����h�dr�1{�+ʎ��"p�KК�c�rE���c�N)�q/�"����I����5�JP���x ��fZ�ҞL���U����)���-]�:�5A��>v��/�n��Ѧ5��j�/m�b�*��������b�b�׃���\�%�ΣP���NK|>�]�s!n���0+a��k�_�Orŧ��U����B8�_���!a�Q����y�s��E��;��@@��b���Ϝ�X�h�4��g!m|�%"٭�ڮ���]��-In;{S�s���I_���<-1GyѰR��p�=�}���7 �|xPX-<ș�=�0X��O�w��\���T�J65,"�'���7Zo�OT�zY�9�0�o�e�k��}�Ӌ�L�KuM�-w�~�jl�)uo��ɔ�R��Iߎ �"Hs��Ch��9M�%����m���^BC�v8<�0�t��)zE�UJ���b�AE���$�m���\S���9����U+��G3c��a.nW�R�����.;:B�6Q	Êv�ZC��Ȅ��6�Ń"�\ u�_��x�Q�{�j���J[_>1�n�`�E̘J�-��~�G���e�<��Z������?�@��1�v���P�����%GP�O^�Q�����@����*o��� 2�i7ड़ȭ���	W�8ࡍ�-��򽵈�s��y����;��1�Zk�����9ho��8��'�����5+$�^kl�r��H�
`�[G:=ph�c�:��s��b6�� �gA=�IdR��_������< ����B��|�^�v��N��wŏ7�b͌�]rA�i.��wMY�?4�b�I�KmU �O�*��;E��pIɘ�1ai�vPcW�zg_�v���H��e$���?��vt/q�vzi>h����(]#=)��JI�6NuZo���VA�vS�)��m3t� �+c�O�/:���-x|P��(D�����U��z�n��p�� ��9C�n���D�4�����_~j����(��}�^6��s�j�!��|��?���r��[B�"~��Fvhk�ɣjm&��\��$bX�_��RM��n�-f�FT�U�R�1c��.[�Y��9X�w>C:T|Ň�p3��*H�lE~��x��@��ӻi�?�_�&��xϒ�װv��B���hUy�Az&�d8�eh˿�{P�j
5n�l�E�a�?����D��\�]NBA���N[��M�ł�nX�}hލZ�k�T'�!�Xn� ��4�_íal	m��b�U��=����,������]0�`g"�{rA����U,��f�+uQHhRB���b�(�Ϩ�bG�3�[��� &"IO��ho����;��W�GFQp
��E���6�{i\�m��o})�A|.J���!�{����� ��
5
7LR�23�T�_�����U�,��#SrAVHQ���J&aA1�����l�`���x��$��� I���:$�Z��5�&N�����+0f!@C���
�]�F���;�	/�,��S��?9)���u�"�����3�B�.3�m��3��2�<�4,�ڸ ��`�@���U�<��[+\�.JՅ���gB�a�A nT)`��Fux�B-R�1�8�"ʕ�\�ʍ����J�Չ�mˋ^'|�%J�%
C��H�N�Tb�3�M1�e3���� �u�?,�v�E�Dq���de.�*p��CU�F�`��cv���]���9����	��ځT�����#}LzR#O��'V��%�s�RQ��Sl�&i��!ɣ��#�K��[����پ�OwN��b�6�Ͽ��F���7O����o<{#,������/"P�6c^���d�9<'9��ˊ��)�}Q
�Bq����L'�����X㞭��b��V)A_�O��R��ݙ�I��&�1Tӧiب�CG)�4�a%�N�X� �U�rAYS�Zj�Щ��lG�`"�Q'4���@C��t�gO���N��@��(���[�];�3�/�9QD����wm��a����7p�+=��G�$��b��m�c`IF�m�T�O��B�엷�_p��k�nv��v�K.劬�����/��Уk{q���7ݶʖ9�Q��h��i��ﲞ8rX�+Dsi���Aԃж�t��vT��;ʔ��He��O���D���7j�1"_+`?#W�D��
�_�f%I\��'� �$�|�����0b�yĎXu��g~C�*���l&l�;�Z}������P�e%Z��{��$bh�K�Cy�@M�/VդES�������	���;4^����%<)��2G��l����,r�hqĚ-�!I$��L�s���r٤?ΜhwR�6�����P@�Zn�p��Hvhb�z��<���%�JHx�v�0a+L�ߍάa��j��ߗ�촎�z�2���g��"8�ͤDT`ѫ�+��u����[��#N��'��z,���[�������X�ҪsɯT���Zk�D�g)�Hn)@����_*�+�bw�����v�/�E`Ti���K#ˠ]��7yk~Q��<	�Y-e��
���V�ǳR��,��\
O�_J-��o^\[��P�SZ�[;0G�eJx�	e��N����a�tS�5�?��� ;x��ٕ3��:�Ӓ�믕{8H�~�R2&>Q�S�0��ќgKx_�=3(������em��j"��XR���Ě�i�Xa�ר�V'��`�bR��rR�����xR���"��Vv���˰1�	&o� �e���5ӽ1E����IaĨ�� �������ȠB��n��d�TM����:+��������ѹV���6�>ރy�'�7��t��X�s��x#��W�˱����W����+kS9r��o�)����q�*�y�+��ݥ?������$�]2|�8?�E	��ƺ��_���6������lvԟ��G}ϑ�w$�q�s8s�C�Ԅ����2�-'�$ߒ��r�&?�53�u�W�Tl��q�7�
�Ye���w�U�ISo��%��;�u��Ư�l�A] _�����b&z�LKez�� ���ofNa�E�$��v�\�q�%�����\����3�~ܐ���$
��\�"#
��}�`�<-�$�5Ɗ}fG��.�ZV<�}�,��������ԇ��'\?i�l{�u�݅[��F�)�"W�Ҷ�II�1n]2��M�T����@�7�X�W��vP�c&Ɔ =�8X7<h�v�Z��Q�<��f�N�2>�OҬ�o�a~�n]_�ā�Z�e��=���{e�a��n�%o���J`�5��I�����Za���J���RҮ��{|m�j�e�Ķ�@�H�f_)�NT�����)p�D�l��;���'갊HC����w�SY[���Y'��|*�Jh1
���!�V���?�������66�'d�54�k�Ų_�Y�w�(i4���|��ՔC[�l���؀�y'|i��H@}�<�	��뇁�k�����!Lhdta��4���7K�k�7vC�R;�V�4�<\���z�GW�	B8�"���m��w�0
�����]�7�t�OG�oU	.�⁰��P�K1b"��~7)�;�A��uMW+ Ի<�0׀��'\�ڊ�fY��Փ���aC#u��ry9�����V V���o���.���+���H�y%.DDv���F$�[E�l��7��n\fGY������ ��AǑ��z7��Ǒ�^���;��#�p�j��"*��
]�)p��p����E�"�?M�ԗ��o�ib:��`��p�d]U�ο����_��#N���|�w�K�t���֦0s��%��Pd]�b�%^ZήS˹i�VC��ʙ�aO��^�ʶ�sЪI�)�h��NK�7���f\�z��TH�4y;�_R�wOng�65"���տ��=��酶
��9��l�U��sKc�f�͇���:(	���5�
�b���/ D֏�f��(�ꯉ"��w�L� j����]h�		bP�'@��vu�o�, H6��:�q��C�1ۊ��o��>x���AJR�Æ�J��f���&���c�Hۃc��(X�ի�o׌�V���9��3����� ����H{��AІ���sT��f��`�2����xp�H�/"�� \b�[HV�1�z�Rb���{�!W���7I~e���b|�lע}K��_�ӛx~Zj���3�I�~�R���l
`�`�.��D*����)��`m"�y�YD&*���{d?tC!��"�Y��И��0�L/�(��ڻQ��L��?�$�8����Pzgˁ�����[��-]{b�ξ�l2�B����fS�*x~m�l�W��(ى�z2�m�ӑ��:S�f8��KT=F���ōu���gSVAu�\�?u��[�jL�eow��Pq��o�˳�p�ދVs�^�"6�SK3'�i)eᕰ��쑔�E�ń	�
���P<&��|��I�m��RO:��ǔa����TG�(l�ܕ����ɴ���]� �o�%�E��U:�����"Q��r@���{�	vĉ%3��B	tg�FiR���W���X;{�=MQΝ�I��T;��V��eC����ٺ�z̲�����59O�ȶV�W[b�ҳ��B���@�:)G���gn�OCDc2��7���'K���A|A3t�{m?/����*���z
;������D��t,�h�]H�b�$���l�gBr�s5[cX�XC����2O�����h��)Ȟ\q�����I F��\�#�~mr5+�6h�$}�����zn�ȕ���|҈�LRi���� �(v��Ӌq=���7�\B�Qo�>ðr�˒?��H���ט�N�5���@A}[��@�"�Jz:���k�Pb����%F '�a
>�řV��}+L��l�Mk�Jľ1��)�6�[[/ӄ ��v�7C0\m���o��#Uܿj��'TZ?���� !OBS�E������6��&�ˤ�+��,�YH�R��s��܆�/0��ۼ�9�^�r����Rq[�]}"����JC�v�|6��&# �q�`[����t5�x��d}��v}� �1`�,n_m%,z���~�WdR«%bl>�1�d>����B<�i��k
<�..�+�o*���ĩ��Hſ\�S3���rz]Ci*���a���hg-���D��2�qt�Y �K��Y"�����2m�"R �:�a]�f� ��<0��GK\p
v�f$!0���Ӝc��7�5<�=���9K|�#��P߮{��|�%.꫌�k�RV��.2�W[(C��'8�2-��,�
T�� E�+��S�LuG8�c]y�3�-��	!�4� ���_�֠߭
�O5�\��(�W?�į����^��M=�0P��:7d�t���ʌ�����?lS�I�O�/��N�t{P��wW�J|���c�w�zMt`G��H�лJt�~��q��0��e�o��&��0�f���S���<�J3�mV/�}�i}HZq��0��1^q#6B�~[%�
�z�t����Oiftݔ�<�vj���x���3ʋo�r��{���SS�uh@���|r�%Xv9c��}`| g��W��}�Z����b<T�����.���PY�ƣ~��KL�=�G\����E�{��[@�������Ҷ[봄$K��I�n�����Ȳ����V��H1/�{Z;�`@<g�hjV�>���s`)?n7�Nm3
�#���h�?5�jYc�*Z��8�(W|-��Q�0R��b�hI0��������{@!�8�?qN��hI���B�E��dކ���T�l�R��8��;�w��-�$�ѥi-��d��p�{���Q�>z,dI�y!�K�������*e��E�IR0�g�lf\�RVv�2��y�v*��I�����}��4�p0ʆ8	�c��k��'�$Q������F��=��c
%�~#�$�mim5�*�^��R����VŜX��؅�������8�;o� n��2仳2L}��
/.�m_SӠU�I��>�����ߌ+�Q�D¸�G��ZG�R��p?����F�&4?s��������J�PN�Lj��{3+���iiP�{fbUf�+�Py��77��,�󜌰��'T��ý�'���j](Zڣ�tN �:�uiya��XaC�=��k�Օ��W]�����iP�e�S��ޫ�Hn?W�2'"��H�zyB7>�!s��g۷a$���Gݰ�m�C��9������uv1q5�chS�ϼQ|���ah�t �2<c�H�6�e�H3M3��ⓧh�w�;���mww�v�� �v]�!7�흂a�wq2� �#ޯ��\v�a��z��y��$�Pm �s	2Jl�x�&��D�27Xݿ���9̗E�e� \_Q�'�cm�%�J+�F��w�T �P�TЈ����Wz�2����������
C��k��S=PG��l.���ZC��(��A/������I=�_�t�ҏ��E�}�]#�~HS�p�x�j���(Z�j§�!���C3��;+L:j�}#[u��	��w�i��������v�q�R��������T����5.�n��i����l��&�^8@����Y��6�٬�M�>�#�R����'o�N̡P���D��V\>���`�����s ՜�}����8��'W�\�g�(�4��{̌�?,~ťؘ	�~�xBV��Z�J:]�����v����`�R�br~�i
v�}���HW�r��r[�6&����5i��^L�5@�u�M������:0%u2�V�<H.e����λ�I���		�4�$zN��9�V�]��\olo���A��9|wE���h"7���_I}7��PݭE� ���`*�[�`�{?����/�j��Z���^I(������=�Lןq� �At�he�Sr\�q�{J[{�53'�P�C�|x��n�*M;�.6��JNp��U)�.�7Ϝq��Y:�B=�����t�CgMl�?�͑K�0�\ �C���灁(��C}���aě�z���� ����}&�)\��1��+�'O�N{��u����[��4�xq�+篱�O�hA�P�w�|P>8�]Nn5F�f@��R�NkB
�wC�|��}�����M���#�5BL��J|����,��g��{�(��
���,a�6�����Q�P@��J5�Qy6ՄA�(l�(� ����Ǎ�9���ra�P,BW�k�� �2��d�9�}"��_z��TA帖�O[�t�M�"�V �����=�5ՍEq	l���������c�<�Ϩ��*��qV�o��v!�u�	۟!F�f��q�E��m�H1@��%�����K�
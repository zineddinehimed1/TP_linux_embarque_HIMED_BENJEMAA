��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�ob<{�����
�k��пL�^0~�{�m	bl$�QmL{�����	�z��P�dO8[(�=�Ye�>�)r��~�e�Y�&�X9GP�3��⛔Ev>0��dW`;;�vE<��y��9�.Oy@�&p�����!Xd���]}E.���-�_�au�,�݃��z��P!�&!"�51�y�lp�*��1·�ݥi\!7;��H�88�~�����Ţ�%�צ�� .�D � %�#�����ڭH���Tzy������*RL%����w��_P��^c�t59_r�S�h:��p=&4Q?M#�>ɖ���vJ��Q�P� ��6XƁ��k�rP(9�����y���(2'�����[��Qw�'�dE�|��>�����s�5N6]�Ï�d�����Ja�����,��4������E[\޻���?��jc9A�3K[�h���ݑ1�[ҼIw޻�Ã��v�8��㚏'�$@к;����Pn�f�yC*��� �t�;��)����z>�<� ��)j�9�vE�#ԟr9w�gv�c�]ܚ�n��([�������D}
0a  ]�T��|:M9Ϩat��r�g��*�����(i[>�QEUK�?~y�������]ڤA��'�✮"�ڑ�B��xK�+�!���`aÀ�X�(Z�Y��a�x�ݴ���c4L#��e@Y�w�v7Kc�S��Q8����fԑU��Y�Ŕ�{z�,��K���|��'����]��v����&V��yz��z�V�u��z�|�R��уĬ�*�-���_Y�K���8��9��,*o��b9��rw�+��]�J6 8�}����X�G�8�ltI�y\s����{�/_�B�-�-j&�!7Jy��S��
�sg7�&	Z�Cp�:��b��:tc�\�?z��wu脽�nA۩�8�a�����:;�+���+�N�Ԉ�3U��u+/�܇fm8�
R���-�M��
�z���䡐L��Ʊ�NA�__��X������Tk̋���mNJ�˺5E�ؖ{��w8|�Ǜ�e�i_\���=B��c@����l\8��xq�߷+0p����$K�ר��̓�@��ǃ�1���NnzSR��ĳ��ID�vi$�  �������t�w�rQ����0��'� ��|	��Hl86��T<ݰv��g��^D$�?���W6U�$��g���C1Y����5�`�O���ÉJq������Q�hY��Vᄑ�<�̙��h>���dƑND擨x�1�8y�6S7Jց ������]	�Z�îݨ��ښ��t����l*�сy���j���f�B,Ϫ��G"?��E|m�FW���ڈZ��4z��G�c�:<)��xt4A���,���3CPu�܁<T��v��gk��B_B��O$<�.�g��M�r�t(i��5�4/�E�T٥q�����+�cLpGE2��p�>-�`�e��Alp�'���N|�*P��0����m&��'c�M�W����U@��0�z��ǐZ�yC�."�0Íz��^`ih>R �x��	�|F Xh*4R�RvK���"�F/����_t�}�OQ�r��m�^��k�x�l���)�c�0���y�m�O�	>d���D<.ؑR�����K~�C
_����g9�g�1��l����ڳ8��ģ1�v�x�Ը�E��c�%_ef5³)�T��7D�%{�ߤ(�Щ�[3�������O��\��;0xn��q7�0���8V���g�!�!��"@��1m��]Y&��`	��E
���ܬ��vҀ|��ꮹ�@7��CĔ���畨j���HH�%<Z�W��3�>Q���>�˺�h7%w�"�	��:��iL9hЅ�G\����f����b＀��5V�^XBT8��2d�{h�<h��ڰ�M�,�k���4ù�b�=�K?��97�����*T8r�h���(�E�٭�a�U(�΢��rTo��/^�����c ���~��T�M�YV+qz�z	f�l����v�����Yc�,�En՗;DP�>��T��*HR�i/o�Tԧ��y�ʡ�
�Ѭ�f���5�V�t$�t#��hE�2���X��|%i��7�`�҃t�(:��8Ri(���k"���ұ3����s�?�[�Z�3#���ٲ��é�_�8��4&��F�Bp�-��&&��GUV��j�Y���xLi6ة$�{�5bgtc�ZO0��3L���~(�ZG���j����W #�gh)D��t4?n�O'�ᤒ 8����=�϶������"�9j��K'���#��Y��v[���S����m��������W��$D�̛����s�\D�U�pQ|TV8�v�>�B����/��@��8�;�7����f�d'��w�3�t��ML%-u2ɳ��,������e_�mH�DKʶ���J��t[���\�C����cr�u\������
����dR��r�N�'��z�&����ȴa����ℒ�7�p�}!zހ)�X
G��SC�:�SP���l���[�k��7]�W?����h�-u��p�����Q���t,ҧ��d�/�F!���&Zfu�/��ܕ{�k> g�XQ���c�x���V��Qd��Q_9�60�ʟ���^�ڥ��VD7&���|��T����<h� Uf�A���P�e�a�0��o4	�,���1�h�]��X�Y��cJ/�$�D�rZK�R��E�{d��*0�hj�8�.9Z܉�"_�Tw`���3Ԭ�����w�K� �Vr�If]�͗�����c�.���Hߕ��#6aD����ȿ��W������_�Y\��%�O��7]Qa��o��3�O߅�Q���1��`n��f����ܾ=���;�UᛚQZ��Q&=�j�E}>�䪺/MR���C^<���,U�S����4��#F��'r{��w��A_�юAV�ξcw�"#��Pe�U��L��o��	�����%=�fZ�5I����O�㘇;?<����9w�o0�F�B'�@G�r`S:�LL��{�ᦟ�X?r]�ٞ[����/�������"�@3���:�����E�%�����/����EzK�r����c<�:����f&�{�*�9&�՞����k�K����O7Bҙl�C%*~�����/�Zl0��N�˧�rfG�[r:)��N
�hd��k�̉�Y���9C2�3e�����Ն��S[-f�P� �w`-���8�a	�{ssP3Ce�h�{j��nD�a�=}���/`���W�2�bP�^nWX(d�-\oG-��f4'o"�^Ƈ�)-:{WK��ӕ�E���UB���G"�$�C��4�
���Êްc=��Z�D���4!�Z����=67��j�M��:�:5�/�K�u�A���Àb�'<�{m�Kr��{��Ӊm.�C<�d����\�֋J�f�_�~Ȳ;:=�_�Dp�	�}ٳDe��,��t:���Y}�{�0b�[��h���R��Z}v�ߌ������_mE:c��˰5O����=�f}h}�y���4@N4]�R6؅�Q�3��Q��c�0I/ �!H�����b���&�������2���{o��4)�X�q>WK�<h�N��*���; 58;���u��}s�t�!H��5sOߡ� �Dstp�.����u���ǶTI&	U��/ä�� �ʓtZ�B�ERePOX�-ɳ=�b� ��3�A�2s��K?	�d�YzTV�&�*�I�Q���F�Y���V�٬cp+�Xsy8��H��X�.*��B�5�S�Q�4�#�cUR��,�� i���|�X��4�A��bV�-�i�}�=�W)�������t�nԼ��X�Y-����
EZ�| �􊹓Bj�@S����<��dCGjn�R|�rqT�0H��w�p0�#��3-z���	�r�O �����K`�9Y��[��&;��"�W�Ë��I4۾�zu�D�0��h����������Msy�� ��O�ˎ �|��^+dЦ�ȩ'�O:�ϴ}�G��c�^��k������y	�r����ǁ%�>�]i��*�l��y|Ά-��Y�/#0�ⶫ	T#sϥe;�c�G�ĳ��{�F{��7�2X�	П�?���Yʓ�'�4 
�i81z�5Aܗ�@w.�ږ���Z?�k�o+Ǐ Y/[
ϯ��$��R����"�S���A�i�gh�\m�%!D� �L#�V(�Y���ꗾ��9|�-�"�0��hqI�y�<<8��#�Cx^?�J3���=���7��
s��r`)�vݐ�>�Z �NC��E]��h����H����`?;�T�54�T �0�}e��] �֕5��Ŏ���qi� l �ȃm�px�	/'�{>��R;��c��!��b�8�����`wӾ	p���"U����W͟РU�Z��_�#�_I1�t-)�.hځ����Jm��)�G�.�j��S�*�Y�q���Y�/�Yy^�!��q�*̫]����3��
��ڑ86<5ܝ,=&��4�� �-@�
��0"��EӸ������w��4dn�:��}�!|y���gzA����Z�ۢ��u�T!}��9�F�WT�T��MJ�˴�A���h�)�8�(Cn�I��\����)��{���`Fu*�%��u���F�-UI��w�Dn�ڛ�.,L�K��[4w�P	6���R�Y�>�����v���P� ~ڤ�[�wI�,FB���|��M�rG��uy>P�
��鿅�����$���_��HԜ�o���Y��x���|�j2�Si,�������&�l��2�=��FjX��W��x"���;����\�(.T��;y���Y��6Ù�OZ��iV]3��f�L��h������
Z?)�p�?�Q�7N1�X�|��$�0Fý8 �l������1�.DZV���a�IW�%τlO؏���&��wѿG��o=��y�����}p$�~9��T�}� d�Ro�.� �������e҈]IN:�2[[y�B{�/��)�{���@O�7Nc�e��g�����%,S��ֿ����u��`�+����
u��Y	�3u
������Dw�Q��G�f]��HX�Ʀǝ�j��DS����"<G��d�˼��	+٧p�d0!ۢu�֣2�=Rq>�r��E$��/����8�i%��}��ɋp���
l͒�)���.k�͵�n��=��]TbY��a�D�X�yW�D���s��d	�\."N�x��'�� dG���h2�;�L&N�G�"����؆�fnrN��p<)�a��Tn���igs����U��(�����ϻt�;�߰��0���`���O�"42��Q�%Vm�ڗVB� r�9 ;��2ن�qP2�Q�?b���n�<��2Oϕ����"y�^u�ލh�OA�t�h�/dS�J��$�բ�;�{�
�)f6 ��#̩^��Ϥ������rqe�@��f�l?8�]����O���𣕯7�M@��6��o���5:��7Em�@3�X=v��Q#�u:e������ڸd 8j����&D��7���F2�xbg]�Ѱ��޷-	����l��qQ<j��Ir���������)X��'[�P#�P�M�:���**))�U���M <l��E�UP�9.b����J�+?'�Z"�9�H�+2V����5J��x�z���8NHZ���"������ �:���v�v(�� �k)�I����Z�<�9��z�5���]��7?��;��3�f�鎇g�w���[���$B&`Q
hkqU��P2�0����|;c���̨b���Ct�q�4��)�(�����n��0(݄�[{o���JtMkֽ9�դج��<�F�����*!e��Z�,Y����;%4���\ϕ�,�!��&��@6�Ҳ��j
=D E<��_t �iC�Ԭ�ͼ�#;�����8�Z�r��.�0g͍��q]y`9��­x��Z`�a*x��|p�a�0��<�=��^�ظ�&����I-�yTt��D�ތ�P�{*�OT�뛩]|ZL�K7��	�B#e	�h��n2/1�Cbm��i���]�-�mi���L�z�Y�ZH�����MO�=�8���Z���J�P��	_�]��S�B�UyO�� 7AE�{�����狳�K�����#ju%������} cV��D٤�I7��/����FG�'NK�<�W3d��xcH�����~�[�aeHB�d�� *0sQֲ �q�3X�i��-.<9�(�����2�Sϯ�o�M��o�"���o�W6[w�в/�2���,v#�R��;P�+vRX�Tv�\�.l��ؑ�`�XXa1c��
8��8��"H�q9T��avT�ll���T�������"�F���Cl;#3-8l|P����`dX����5���\�D�f��<�T	 ylg��.x�t��nCNI��&M��e[���"�le�@��@Zna��Ph,JSEKL�>{�ʠ�%�p�
8	� Rq�ݐd�^�e�;^�b�K���j�Fb~hЙ����Y�[8u����P���\�vL�=�9[���k��0HZ�M7��t�("PZ����n�斲[m�`�F�_�|Պ /�։�@�,��p�#ov�ԶLl�p#�E��=x�N$�?O+��P��6m?�r6Qͽ��7rL�K���y�o(P�R��lR(o��G��$�g�9˄��Aľ{t;ʤK�#��X�0@@uCP��1^"�|-�4x�n��=�ސV�ե��T%4U󞗔Aa�ޘ�7@�enA�9�[):ܑ_|��Q�W8�u&��YĳD��eӲ�Xe0����5Ug|�-���<,'+(�+��Nx ��34̎��vI-ڝnV1��Nm�^`�����|�a�m���Zrڠ��&��%�c�{EX��5�����7˺|�>-W-�62ל�1]p�E}�0%SǛQ�٢�Ӿ+������0y.;;��"�уK��IN�������4"����r�dHi@�^1�I�+���H���X>�bt���lqZ8u̪��ZA��?tT��Ǜ��٢�}E�k����&��$�:F�^l��U���Ы�'��>��D�>�}.p��h��>���<a�[��TìȢ��u�J]ƚ�K��PIaca2���So��)cT"��5�ik+�$�&+��A�;�4<����?�婋�
k��"�{�CZ|��i�{r����C"Y0{����o�s�)�-�=(�]�D�1���(�٧�@�����CP�npp��#��� |6L�E�-hF�q�9UM��� %v����?��y��?�wZ[��Վ���` ��$��3c|�KN��[5�J.�;(�kK9Tpf���!l�"���4X�oS�Sb�z]Ĺ��V������<�'ҵ�Ɋx��?��f�e|�1Ыd;`<[QՎ,`!�̒m/j��]*��2�B!&u��]ȅ�ݫ :&[��|����Z���-��`WTV���Y�yhi�1�b_��I{�软=]�$Æ�+�Q"��s3��S����4�3�J_��#!����2\�8��d�?�!���kxb=z��7��`d��k���l�f�6i-/�ƌ�G)&��Da��I�n�j�Ӹ��I���p+�<{9��<� *�|�%��0`�x�[?��+i�*HA�;]���a�#�pE��G�E�v����ޔG�:�3p��'�{����M�5�:Ï89��z3h&�۽M����E�]�K��cr�|�B��C�D�j4�]ߴz%�B+�4�n�u-\�cj����i�k�9�*�N�hh���Q�n��O�������QU���$�Fic�ш�V�zX0��h���Nxe���&�}�i��3�u�>��4�[AH��K�*��l�������naį�;�!��E�-�E`���z����;t	p�7���j�B⽃L��z��u�H*k��?��E:����x�o���L��x��Ӑ���6e�|�D̥ �)�+�]�����ɹ��kqE�{N4���;`٘`jsJ����F%��;�qf�Oȩ�,��%O6+� ^����;��]>�	�C5��h��I����w0��}iJv�>9³��6����$ܷ��o���j��3�|���%�*�75h�}F�|���%�k�I�D�8ѽ�_�B�T�FOC����,qcgP�ܱ ��n2�t��P{���8��b[q�4��0�9�����z}�w��M��_�쫓&�7�D���9Y��J���#T镻��}e�P���� ��p��/�F�:��8G!8����#��s���_1m���VP�m��!&D]�k�K�d��vp�i��(gFB�_9����N��� 8~*����g��R��ܚ��g�ߛj��;1���sm0hpM���l�yO�/���6(��Gd���/ba�N������Rx������g��NSQ��}�����4��<q�}��`�nY'X���<�d�:p3 �pG�_�x@l��*�[M�]�F��?����V�����@W9��wU93U��"���pN�tJ�sh�����۞�Q�	�'�|��B�,C L��P��X��E��)���FQȏd:1����?�o9>����/� �Z���Ը���M��1qHE�
�M@<<`�@�������L")5t���0E���PύG�6�鄳��kD4�%;b��
267!R3Ռ���j�sX�V�5��c�2��5J!��+��!�gV^�af�X�¸(z�|�[�����`�[�i}��þة��}��[���˻������˧�P�E���l՝=,�=��J4�H��Ǻ۵ܴK-���k�P��Ȃ���:� �2#��o�d4�@.h�}�W����� Hx%+�d�,�3��!d<� ���\�
���� ���]Q��!��z�4l�IP�h������n���k��F&�f�V��@iw[� i�>)ZDطbf�IAag�۲ܛ�;x$�,��X��dqMKb�����~B�U⟞kqe	i_zsU�<M�%{� �:r��]V�W�b�Ul���G�&c6��=3����ԟ�@�G�n�b#��&p�n����n���'� @]?3�^��0�@� �t)+�%>�3h���*�<l�r,uw�_���k��Y�[*�=Lk�BS�w�����<%�n�04dI�f���e�Sdլ�Eo����ؙ�Q���L��9�
�S�-ڜ�����IMǼVў�]�Bōe?3�_��-'`�$����w�������^���2{�z��9;\����Ŋ���v	e"��Ū�%��U��.l*(���MA]ָ�	djX�c<�L#;_)�%U�u����^b5y��������U6�D�1#���xQVv���g;�����hK?RŸ4�h��?���[�"�9��'n̖�j�w�S I���B�z�G��}43J�:�l�=���HI���}�t����b�}�zE8�dU)"�-^-Q�`����쯒Oi�����/�;��'�Hi)���!?`�8X��dDj+��=.pѻ�*C��;de1���|��@��p�C��gSj�z6�As���%���N��-���8��{���<���:�3�Ǩ�3:�� Х�
Y�� �3��*cX���Ş2XDŀ�.-��r&�W�e���~����=y���Y��7��u�7�$��Jv����JYHF��I~L�a���dm|����:H@���	`Pm�[�2A�qI�=����R�32��R�*��/*7���H_J�C���<�ơ�D���V��س��=�(}ݯݔڴ�Vvz7������N+Eo(_���\!<ע�X̰衈K.�z�T�\H�f4�)IZ��'��K���uT��Kh3} LZIc\?�m�K'� �r������ �e`��7j䆦(rP��SY�\����p���;r�^-}=N�
cZ���kĘ�>�@��Ubؿ��Pco�^�:v���͑�u��x�#�"RS8_����L2�ւ��M85�R�0q�[��ą�1�0�ʥR�1X�Z1C]�4-Ԑ8�(��2]Z�H��o�G�<��5�=ψi�zy�i�Fp}��%�����\%�~^�~Yh�8Q���4C����/�����Y�sH�)��;@U�F� ����]-NW�a.e�&���$3�[���b)��AY��	��yy��{
��=Q2�L�|�&`������|�[���vl��g A�C��2:��R%'և�^�Ɠb���&��O;:��M�cy(��IPS5��r�wG��4;�X�X�&5/�h�H&�"}��'g��ܤ�WYͶ�'�s�1����mhQq���������6��0�<Ԧt�zT��f��kv4��
b���/��0r:�b�Ѱ+DoIVO������7qa�㴉��(	�1 �0*��\����N�Eh�U�ui�	#���{^�M�an��������d�3v�z���g��s92>��S��r�`�U5��ݮ<������að���X��=v�m�����z�98]󛦧p�S�t+J<ie$��`ښ�f�nz58�Vc��!�i;���971��2`	p��3tu����/d��}bp������Ʉ��@$^Й'�â���e��L��M�?��(�b�L�]b>�ךD-Lp$��_���O��?��[�^��K
{|/B���XW̩0*���ӧu�`fp����Pc{}��z�g-��@W��֣�;"o�������ql >Z����r���1,�e.�ӃY�+�������ƌ=lݠ=�I��S�	22���Xt�H����� ye��7*���E	��9e�\�5���*wo��#����O$�)5(?pȬ^�]J�vEe��I����ߔ��m��n�J,��}n:9HF��aG��.���z]N�͎l�/��OR���=A�~u�Z�8���RD�򳞉ѭ��Z�`yIT2��3tfc=u<�?�y�W����R����M�jFP���}//kg���6̐��=&	.�I���^���LϺ��� �CJ�Dآ2K33�x�f�p��}���h{��������H�-_}�!��>�������fg�%c�q_
�xM�?>�޸�5�E���]	}ֿ޼��� c�6�y��;
�`q�S��dS,�ZO��>�Ү8�c����Sp�ܕ��G_%Ihޱ�ެ@�?:W����J���q�I �|����^�YH����홍9�@�UR���N�a�{g (xI!WD�>F-� 	�5sK����A�A��ʔ	�jC���ۮ���5���q
��z���KL���V���.�e9�S��ê�g�磦vg�؎4�h�:���,(6h#I|��Ձ��]o�r�mt-�m3Lԁ���Mx�6MS*�)��Zh��"X�ڸݝA
M�5qvVk2<���2+������w>/n�Gm��^̻�Z�=u�w�F��Q���OӢ�'{���w���T���>��7���k�ennp���I�E1�GK��y,?xS]%O��O �ġbE�B�u�~����������V��V萤��HM�	ފ+��=s��I��U`(��݇3�6��<��C����.	@��KM�'@�W�b�D�tk*��98#fM":�y�,뀂��7N��&�".=tꗭ���r$o2!�A}tz\��a��Q���[�2r���jF�v:ȉ��e8�{�@ l���k@f�vI���ť�J�M'l^<H5L�Ǹ�f	�I�4y�-2�8���e1D\��z�h��b�x�g�wz#=cykK o�'���Y\���iA�C�#4/�s�ؔ�����4`~��8j�ˀ*>A��&�oH
���&2D�eɿz!�11�f`������^6��Ԉ�1�ư���wU3������Z�1�;R�/���K3K΃5N�߀7#�7�tLVā�P��X��묮���$U��!p0�u#U�����8,�0uD�3�	��W�Z6����e��.�7����ϲ{@O��6�Hv��G"v4�e�̙��%�4��Cֶ�9p��
��q��k��W�a��r�6���M���}�4�S�//My�-J��Z�S������7�W����C<2�i�>7�zY�������e�GS��!,��י��T����qJʰ�~��·o.^�V+�R >x��ӹ����ş�y嵂}�vҼ���|���im�w������s�w	�Y' `*)��H�p��+�ʜ>u����|D���sV��ɏ,�}���J���f*��JX���ҲBV6F-�F�8���2���|=6(�AP���1�r $�ݾ�.��WZ�G���{�j�F��L�|=����R���q����S��[�U�D6��!�A�Wth)N��QB��N���	��O�)c/ֽ�"��F(QpW�.a9:$%��/�mB-��YŚ&���T`Fq�NY7L�����T��Dpu��!g �c��w��:n�F
)͡��Cq�� �F}N�q4����RȞ8��>&h�$�?G��1��1%6hF��HM/��m\�,#*�g=�>��ke�C������dM����F6���eڳ��b@W��8d�F���[���щQE:���qc̟P���@�}{�R�@��,
P�z="�+��z�74����W�:;���z�Ub	�2 �H=����h;�d�.?RD�g�o_Z�};h��"ijOVp���^��	� =�+��LV_��҄���̞Q�
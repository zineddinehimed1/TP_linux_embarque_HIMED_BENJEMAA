��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�i����)!��2�3�Yp���4��ø�����;����g��~�u�a��A��L���I c�N�5�������54�Ѫ�E��́C�i6��X�0R�SmEW�3��m��̤�#"�N��@�����b��aL��O݌2%f�E����t8(���~��t�;��5���ޟhd�-�9�d�/�lA`��kɔ��]c�jx�)%W�?�Gq2��e�u�F�z�=������h\lw�\̑��5��e%��3�����-��7������õ�|�ᒯ12�V�]�b��c���%$�m�����co�c���'�x�@�P����O�->� 9��ڛA��][|��d�D�3x.��;ш{LÝ'[+��W��Ak����ZMyM��	Oj�Gc�`�.��8[�n�f̧�/�N��f7�G��i�t�X�|�z��U�:�>]9O��W� \wN�S0�����6���G�v\��x
�?��eO-!u��|*�00� �AKD�)ŒJ���B��!���z8WU��(��d���W{ηא�-���n��y�}5~�WM���[Hc�*4���7=�E������/e���ΰ�\B�n�9h�)��s�~3
yn�H#������M,$G�u��ut�A�ak�Y|�b3�m�w��Xu �9~ԛ���\ײ�� �wQ����E���6�!{��! �r")�A��q6<FЭ+8��f�}ƫ,v�����I�2U�����as�#�?]O�k>K�+q������_����� �A�_�x��� z4¿-"��-^�DϿ�Kb�y�ms��rG�d*F�@��F���n��2��$��UK*�6�w��*�0bP-&Qo������*���K���Fn�\����C����U<Jy^�~��X�WҘ�j���
������[l}Q�@ELWd�(+%��9[@@�3Lh|�m�Ջ����Ml�b�s����.��b�}\́g�ޢ���@�T&r7w`�+�������t��y1[���}�b ���X���Wfʴ���Y5Φ��r�w=T 	{Ah��01}��k�3/Cc^,��z�?epU�����-Wq�^��o���$�b�����V����I������w$a���?���+����i�SJ��p��M��>3EݒpU��H�s��^�b��tf�4t &�ߤ �� �����e����ժ�_w�	sj�Ht�Hť��2s��^���H��iI��Z���qF5 y
}n6�W:�|9ݸ���+�%�K����|�{��o�����PB#r-�Bu�|��M�����Lמ�X�w�Q�W�4�������y�F��:�J�؍~)ax�e�q�8�5y��������;嶀��^�b����'I+	���d�<�ܽ@�����= ����N*y:�Y.���E��ީ��>��U��7ߵ��j�x��r=>�]��}h}�XQ�sg��׭�ʨ�L9����_�m2���q�*�{��9��0 XaP�����FØ�a4�Y�:�)t��|����f�>>��}��E��#8�[|���̬V"�|;�]�O�ɜN�<�`���{�Y@R��� �Y�'��v)Dac�nG��=��aB��_*Y��8;����t��M'֏W�5��~���&NﬣP91� \����pHB�~м,�%��2վ��a�VNm���e#��W�yZ��뒅���B����\��:i	ޅ���V1���(|�҆����S��\:?��9ހ���lv���`hEIdN���u[f���͹.��~i=�c=#qGz��@�M"�X����ƤF��3S{_�ų��2��Ӝu�Nu���9����{�b{,HNS�p�j7$������=�b:�pEBN���7��"�Į8		r�W�Bf����gȏ�E̛�_�E�"N�n|9$��U��B�G�#���Y�4��[���-�*uj��,��@[�4��
*g�Ԍm�E�ǝ)���:��*yh�ˆߎc%b�k�J��j1�
Q?��Q'�|�C2[]�JI#�\�<�4č�p������C~m��'W���uo�PD�\Ƒbĺ�����Z�	C���4��;���	����u�}��	W�B/�P�o�TF�9��wD� [�~�=t�%;�P��0�Lq]8�[rD@ۇ�[Q=/h��jv���8_�oH;<I���d���y�)7�H�{	"���pj�FI�9����M��^z7 ��=� !�ɳ�亵߻�[nZ�[ǥx���"����[�ńbZ�BQ���Rۼ�=�l�*�XQ;��7�,�o<�9؃��_$�i$T�M}�,-�����3�O>cl1T�;}������Z�-<Q/�{o�mkɰ� ����K�ǌa:�F!�2s���&�Ɲ��b�cL��c@b7��W�\�*���f
4�-D,�� �v�A�	�3=D��� j?T�`�>X����@�cm�UD�D���K�u(nwY���*��;�u�zcl������m�u���
�iDb�[��e�����#�n��a��Nsei#����_;lr���[��Fa���$�_������g
I	7����}7ȥ���6��?g|Z���h,q�ރ-������ CW?���MD0�s
������?�Xh3QR۱p�(��(u\f�7F'�w��}a���#���=�M�>�;Y!�=��a&Ϩ#@�HU+]���ѵ[��͢gY�ԥ�/�C4�k��Eʢ{��b A����М:����AR��ƨ	��"�r�Ո�Ǯ��8%9*�V�I��D���֥v��gm��pqs�����ߕ�>�7Q�wxE���<&��g"E���u��T�`>OF����vfh&��wuQ!O&��xn����X��z�=n~\n�Ufk1����j�F�:��t@}��Gn���Ce)XJ�\>Y��!�)0�졨�}&$���iqzw��if��E�g��	x��M1=��v���X^29�ɲ����7��㈤y#Ⳡ���1�.g�t�҅��D�o'����Z�pU	����#(��ac���� {��w倰�eZ�R���A�1�J���ZtZR�ç��,���OnNb1,�?��2�����TWyF��uN�af���KK�d�x@�\���u�bl㼒��ULr���sN��M�n<&�`ywbB�;Q��� ��*$�N2���� �ai�� �Ue�WRK���� 'A����_G�Q,x�
�N����򄗝�Vfr��/���̝�n�
��±7��=���kt�cD����ݔ�Ϧ�P���IKޅ\��=�Wu��`Li*鲭�����_H�������|����#�!��6 
w��/ٴ?}��#�c�Bu؈TBM�{$:`�9R�c!�D� Z{=�m ���SH�=�E���[��[F�o��n�uEg�Z�̦R�}@�=}s0�qC��l��,��lH�%IVC�%qE�,!zj2J؊���79��#EG���}|}��SfU�j[ S==���!�AӢf#2C�8��f�Ɋ���?�_���{l{��L7�o�v�6?31��U�)�Ө��DT�SHP���[��0��;��Hr��>�Q�@l�*�!aȶ`�J"�d;"x�������`��1��v=�<�
y��I�Y�#(,���?��
�l�a�#�#�4�p�aK��5{h�p և$\:��&t��P�k sp��j�>Z���}x��a|FuH�GR��1{q�Ag3�B%���̤�\m{kAi�� �\��4.����ƣ����f��}^ESu�VS �/ ������L�����bzl��"
"��"�?�Cŏ3����K�����#�U�W�G����2�/��p_�	Mo�E�mB��<�t;]��}�["浼�����0b��0��]|+��1VT�9dU�	΄��ybc�A�ֳ��YjƣTik�b��I�M2�\}�d�D����E
������ ����~Jw4q�V�,�u�T�Qh�/�k�7���\���/�Q�S8R�P"���k�E�I�>㌿�|�-]�m�w*0�z�Ht-���P��݇l�[�O��`�|i�7#������5��}��xD��Sk���h<�EKL��b��(~�<|rQ;m��?��x9w9�"� g�'��Y*�J�^��Թ�:�.��jD��f ;�`*ۨ��D
�O�R�V2��wq�z�,�z��5�8=ԭ��#ի��7��_0��L�N��a8�E�[H�m�Y�*�N#�8������[�G���g>�Eٟ���D��π�����*����q7�oU�����q��-�U�/o�8u�ȝF�_��K��W�όͲ;�����%�p��PS�E�)!��2�
���Y�ky�_�Z�8j`���q�ي?)�Ox����7=L\>��&����ц���5e��ҕ��<{�A��gآ�@z۵�T}0�Uϸ���b��Q����z�~Q��2��.4�Z��_?5�B7)̟�$z�*D�5�P�l��c�X��a�tg��=�Q]Rc�yU�8�
c�K�u�M۵�:	̀D�Ԩ���r
�
�c����&�����g
l�:�[+IgCr6b^��V<Zʄ��6z���Q�R��Z�|<���@J�Z{���R��ƥ*"/�N�W�]j��]I-RLY���I�9��{Z�q+ߍm&W]�[�J�a�>�A�l�\cB�@јL��qE;�,�V�����X�#Z\��^����>|A<��s��Z}������*���Yy�D�g1���Z�$����͒H������J�o�
�Yiu�um�&J�����YU�q�U�" Eka��nc���tJ�8�@�2�r<v(�6kj���>�;�m��IsXo�����4�-4�~������|�ǣ��[a�D,���'bX@{��Қ��f�&�
YK��w*�=���[��R� �>��׭�`�����orc���¡VK �������9F������l���n��~��P���Fuv2����dO~��!�J"pڴR&��y�%���g7�ג^��\��=�֤r`�F��B]�v�>:U�БԀ�b݅��_���ӻ:����m�-2`��kx�|��WUY9� ��V(��E��Xbw�f�m~Bɷ?�n��_���V�K=��g���/u���<�^jĳ-����P�Y�P'c�V��G�f�)?߇���?�MC	�����
�W'E�</{�"���0�cQ��:]6��	૕r'@PG�v>�Hq�U��#z�̝��������M8,2���!F����?Xd�@b2P|w.^�c>�g!E�ar�S�k)"%H��*g$AQ�H���!�!m��^�0�v�I
��K��j2LC5F<����W.��DӸ���ҝ��ny�������8Ӟ���8a�Q�w}�|%cR�����	�8�Ed/w'�]X���|��K)$�j��ۊM��V�rP�Y5��:���`z�'����p���
�C��a��۫�Ι��1ԵJ]>&����;��@Ef:�2b�<GG��� ��C�Q��9m}6�[`�$�}+P��4+��x1 !�77�c��3�c4�- ����[c��zO�c�Ei�Z��q��i��L�扚���h�H��G���ؠ���	���*�q8���l%��ov~�J����6�<����K_�+�6�����+ۘ�[�ހ����Ͳ��x��φ�܃c^�R�k�^��qS��d�o���s���zɔ4��&�,��P�N�y�S�{�$?k/��i�_��䬧��V�j����l�W)�-�����o�����gi!�	�� ����붸���"��vk�]���E)`W_��Յa�^;&e!���dR#�:G!YC���M��
O=K���s��h��;{H��ErLw��TÆ��^σ���e5/�>�%�Xz&�n���s �D$6����9G?�'F�x��1Pyg�F�,�5��mMt'E�l����@�k��,=\Gǳ��4��Y�Zb�����3��pѨd5�V�aJ7��7iT�_�2@{'m�ę���l�n�5��x�c��o��d��O<!])^�x`D�~ z��S7�}�ho�4����o��.�iUy5	��N�`�T�>p��&<���NBlGo�W��%�Y_ۦ=�mn#۽���pi^����a�>��hO�����J�		>"|}6�"��D��k��2!�����9��b켪J2۱q|'��#*�O.�({O�^kxht�����+���E�&����~�C_WP�쁰o��g�����\%�G��D�ґ��X�n9G�Z���n!H�M}2��5|�`����kG�s�unn9���e���v@Tj�T�QJn%J&w�
;퍮�=��7C�-B�y���^�~c*I$lfZ�3���W��A7�7D�a���X�PPj���#V�n��Ժb����*�h��������ve�����J-B�|	�\t?�� �Z��U�����Cb��}l���dWbe"�p/?���ؖ�Oz��iq��1��	Fm���>w��-����o]ݸ#��k]a�{6����*�O����f]��ۮ�]qj��!�ꮲ)ZVV��5���.C!lj ˏ�K3X�"JUv�p���C2�8�,��]��D��;(y)O�^��;�F44D�qq��H��]}�q�����8������w;���Q8�J�x_нv :!My�=�S9��w�����3q�%��y��2%�g��� �|�*�h�t�Z��5Sx.�~|M��f���"���d֡�c��1�T���L�C�s� �_4_��P���i/R�)^��#pix���zk_p�a:�,� !��P��_uB�X'�b Ӝ?��
�g�\����$N��O�95��Si�9q:I�!m�a #����O��g�k
��=�B�s�,��P�rt=Wʛ+0�y���3p	B��s���_g�����X8w��&��B����x��'��9.����/��ן8�y��&6h�:0��I��e�V"wHf�S��������ɰܠ;�������7�j]Fx[Pa����`��9�ݡ�u�({1�Z�7ŋ?Q�P� ��s�.�-�@�kו,5���Z�5$i���gu��hz=K3?�s������
���1q(D�(P�h~��pj/�2:�퉲%�]�+߷AIe>Xw��D_�`v[�������p�{p�`��39�]j���H��8�sD}��C�_��_����]�-��'۹Nb���� %(\�Y�+_ug�:�k�b��AQ͑�Eu+�7�w6�8�m�֍m��7��������mYgW�B��&m�� ��Y��`��<-���~����
!�T#�!�H��*5LzS��m�CR#�=�G��7��nVF�w����?�#�)��D6���I�tdaΐ�H'�YN+�����(��e�P/�]��N:{�3cټ[�k@�U ����on-!h٧w�&gf�)�OHD�0Y��7C���"i��A$�@��mf�ʩ�=#;6�\�d&���p��ښ H���D���m�I��Jkކ�x�@ޅl|	�k��7g꣼~��y[�JL�(YBL2S�ɗ��ow
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2ic6�Y�FԜ��m�V�FҲ5�X_<��V�eB&(�=]��C���~3rM�S�W��ʀ2���lL�
��9�eɻ5A�ڶ��j�)�����@L��@��УDd=���t�e?J`H�PXװ|Q秐FV�-Bڂ�̭ӧ��Y@��~h���5Iα���8��1 �;t�:��c����߇8��؅��Q�)��c.`�\w���~w�9��Ub;��/�֚(g�f��/�E�o����Tֳ4E���G��S��>��� �!,'��c3j�'�݋��&�g2�����mS�ؤv�{���P���mg�;��?H��:|�Q����A_[N�e_���')s!�#T�E:����ɲI买ђTM[�ܟ�9�DoWl�i��dN�heq�� �4 ��EO��F�[�j^i"��"qUǱ�]=��i��B\��m��=�9��D�{Q��1x>`��#�X�� ʎ�{=M�_pJۤ��l%8?�CO$�g1�q�-�J�����8FEu�HK��n��娫��P�kY�`���{��n�;i�-J�jb��Vu�f4�!�LN���P�n���SĎ�}�B���7��|]�Y,�/�%��Z�^-� >Y}Lޑ&��>�����R�����%�0g!7j������3 �P�΁�*p�(�W���y�v���(4���v�?�o�3�M��$�p�W���8X���35��z�@��b��,�S�]���m�Z+��-��L�~�)��P����.	��⎿���ґ8�j���¬3,�������Ҁq�í�;���^m���lm��0d�`��8�� ��
�`����Y��Q_Ny�&�2�/�L��к�ȴ����U}��0XzE���Hy�'^�U�2A2��G��{�5`�8o_!�~&�QI��4c˺�0�y��ش�Z�!�2���J���0�Z	�܏F�z��2>���K!I ���{�gr��ڟ�m:�5Y@<��o8�Ž��l�����\m��S�_.OA�~)�ݔB!�@1Q��
��XN�1����WŢvS�vƶ���c*&߯׸��nn)�Sm��E%}K�L��b>=�I�b�� ���s��j��
-���ށZ�>�ߞ���_����͢��6ǇK�f\���A��3G�F~I�+"%�n������zC;�+@'��]���F*yv�#չ�֣���\I;/����W�$#)���@��Z�҂��
��e� �Kc��}�x�9��(�X��c�;��KTʖ�#�Ԑ��*R4E��V�,��r�v�l���	Ol`Et9�s������V���fc�s��`R��f���b '���^;��P���b �����Ɯ�U$2#��yK(��j��O�Q7 S..b2�^E���������)	�"}�k4[�Tuj[�qZar1g�Q#U7n����`$#Vp�	����5!Ì�M
�\����؃�b�Q�W�X&�*[4<x4c�}��*�3�YX��k!,�4I��ܾ��4*�r���@�e���B�&��=�ڷO]����'�
6G4��m��uP��Hw1�Ws��z���$���!��������K8�LN��G�dRN��@h���evѬ�Im歲#�5�1��R�ڈ���K�t@�'<-�ki'��$��J��'w���G?�� ���k���c���X�uS�T��rT��c�eQ��� �O�g�m�BI2��Iz��m؄.��	p��o�5���<_z~b:���$u^��W}���4ʁ�Ykf�rh����TX�fH���kQl/+�:	�����ா���z�֬]��x��m�T��Iee��~e�ۺn�*ͭ�<��@�A�r�����jK$rU������iL�:�@5���Vf��(�*U5� �O���1�H�����!�F�eDbϫ�g-Kuj@�
A8��
>4J���}�IǙ���/�p�)�d�t�xl>+j��W�ܗ+���B�o|9m��tY��%`purV2˾��db��<G���+))Qؓ�X�]�� ��R���a�Ϩ��t��������X�Zb5%�L�3d�Ӟ-��9�8�)#�spv[IZ��
w����̮�h"�ԺI�T/}���4{3��ڤ{����O*�/�TU��tt7��S�☹��~&�?�D!|d�d���۱�RY�,����u��Јqؕx�$�aS|�:{o\N�-�^%��U��*>���`�����4*b{�7�� J�7^{_�
A���@�~�+3N��A�.�od/��/��a=�\���9W�6������x3ğP��G��e� y�����L��E]Ms&f��pJ��C�^~�a�z�0}X��Ђ��AǵO'�b�D�r	�wB+�7�����8;�>p��?H��ār�Ja}Z��o�Z�	g�֢���B��i����gh�jC �eU.t-�L���g�2s�P��kh�9=��B�V�Q�%���=��_!��]��ɂ�}��5ZۯiG��cf�ܰT�ǖ����]��-��p�x�����̤��o(>c�J�p���/y�5��)=��27�;��L��Q��؊���u=G�� /L��	y~WPw�\�����LƷ��� �5��}�v��L<�q�%lp�=�t�k\�9$%�lD�b���������	��;��ܠaƿ�UX�)�V��V�q��]V|F�ŧԠp:l�Y�KHYS��ù�Th�eb�ZJ_�wAmݱ�[������!!������c�����V�q�����'�	�BB�=n%�]d�L�ʊ��M�{򧳡�����dMr��dq2�BS����o ݙ�5�|N��@�v��|�q��D9���v}���(hOi����nB���_�nF�Uq�+N[n˩����!�E�7�I��F��4A�9e�q�r2�$$�\ԍ2�&��o��ԅ�vc��;�fM��h1�pMw�6�v4���p;�2˰��m���TW1����h�>.AfF�(�*��EW��4��e܊�����6�FX7�ـ&�ʝ�i��ɀ�;P��Ƚ���t]I�D�H�I�A���~�|��;������0���U��d ���붴��}#�����|�a�}+\ԫeǍ	%� dө�Ei��o 3�{��5s�΃ݹH~r���,>����ҝ3�q����ݑ�Ev���\Ѿs厸*t��mBc8�ujrMZD!��=�->�;XV�Ȅ�� 0|�j�~��N���JxnE��Jk̆#�@
H8#2�'��w�S�N1�;�L�Y������~�r���������O<Ex�YNJW�@��"��'��G헔>uHC�4@4��`k<|oC�V�������(T��P���!x��-�=�BІ��|�ϛKѺg�X�`p$#ٙ��L)�����#9A�z�K�k˞\�e��
iޠ'�$T�DO�ΐ1�G̙mE�=���$�Šc�ae��~�Z�6;�۱��{*v��f8����|ӯ_��A�rT��	�轵���ϨR5����h�h{, y�`j���d��À��mE�
R�t&ۆ!(E#5��O�`��]���PƦWD���ּ��w��j�c2?��#�Z�.�fMVq��kM�0�{�}o���;��7��d�S/�;{�O��X-���+�����J�h�9̍9��8zj���k|�|j'�U\�����EbX�I����X��o]?o0ٌ�2aeu�}q(�_����A��+~ύ`�!�*�7-���F�-S�vk���x��j'���6���p&t]hѐ䟠(��(V�ܗ��a�,Y��_�dL)�w��Wۍ�U�z��'MNH\�:��1�����eФ�8�c6�"���*��J����Cn\X�\x��|ql���a�hAֶ��O��<x�y�.��a��-Zc@�D�������/�>��,�t��bO����TT����c�
�{���3�\
�Gj���n��%��-ޝl,cį-<�I]�4��xj�4�����֐(�,�D����^\xF<��M����5�qb���
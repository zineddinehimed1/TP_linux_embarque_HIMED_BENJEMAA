��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"��N3���lAs��7���I��\�d��K��l���}��
��9��z���~��&��-���I[3z�%� �Y�{F�3�6��QF�, a�L\�=u ��@vw��9�%&��H�q�\f�S콎�*�caX��U_�.���eK1-}��7�N���A	���7?�c�0/��~���f'�2��#UX�1	�7��W6�Kl�t���ܟl�b�~�}���Z叢#�o���}�;4���T�'d�x�Co
A����6����� Ot�NC�:R��E o1E���f���>Y�K?��T{�V���m��2kj'�\L(fI�O�?R��U�M�c�,�ի!J��.@~Ik3i볕}+(�N-��)��u�|�Iu��dX�\j����.�ʃ��&i���4�yI�ߥ�m�g���رL�$:W˒�cHxfLƤ���>O,_�p��n�N�IL�Cc9�k�j4�V����2̍M�x���6��<��W4t'�<$&���H-�`(�#�E�Wtv�������OE,���Y��_��*I~|�^�2����%��]��9(u��'0up�*S��*�IM񔊒�(��_���@+a�ܲ_-���l�8���@ϐ�b2�J�K�@/��w�������� C�#Jy��PtѮZϕ�Є���K�ｫ�w��6���A)[�9D������r�az~��ܦ�I��.1�H^�2	sb�����N���>��R�je�9�T���!i�.�eV�a�
��x�zxz ��yW�i�u)Ud��z��Eŷy'�}���]����	^hw{J�x���'�9"�� ?��A�~��a�R�S��0�C
�]�Qf�ν~6���T�0�/lguv�
�":U'�UR��>�+�>�=�\�`U�WU%���H8{��s߇�	?&3
m	����`��	�8o�����S�L�e�����3j�/[�<�	�X\�����-�]�ֻ���L	kW}�T�hb�M��^S�F^� "�T����h7��*��%Ƭ���n�w��&9!o�$?��ۛUۧ��T�u|78c�z����3u���U��Uߎ�&%b��7�OE�_�?��%����vg��H&����J��"#����>%���7�S^�5�6�]�ȏ
�4� ���i�aPMnC�	d�>R��� qNp��Ւ	Z�� ��o��p��*�璉�XK�x��H���ϻL�:dz`�8�2(�=8��&��&�)�<=v��u򈚨�+�����"	���,�A�ݖ_���C�%w�U�t%�X� {��8�5�y~�=���I�ͣ͞���^6Id������Y	���X��/�G���_�w�6�A�A�ຯ����ڪ�B��'�)�.�*�|ȩ���/�Փ��G����$}���datx���C�4�G���hy�F���	�z*��t*C��$�ɺ��/5@(]=�:���u$0*�"HP̏i8 b����Ϥ[2q���P��WPuzNQ�j��E��ta���%�İ����X�p��8��5x�C���"ɽ�M�߃#�N���sk�42&`~c�|�gzF� m��N��ʊ�5�%��D��{W����){���a�	��X��#b�FCr�Ý�=�(��B��%���	�z��i���{i�s�ƾ�o� ����%Ti;�f�2�-���|��Q�	ˇl82'�po�!=9��1�(<��R ZH�$"�B�ˈ�n�����:3c��{�X� �.#�^��êWH´�π���,�īiE𳋊�qme���o�z� ��G==�N�-�B�OF�<t4�Ӡ���O�n��'�]�RU�|�CX�Z��M}�B-��4t&s����.�`k���
۶�E����G�jѴ�i���܁�u��?%���I����2u���]£f['�&��a`!�� ��:g=W�&��������oE����Pm���Ð
�}�'@��]t�6q�R)�V;Z@������+Ā5��Zt���O&a���òW��*R�b�
��e�������b�S����rk|ի�kL�AELWF�a�ݷ���J2hp"�6
VI�;���}��}d��!�����P�6pC\b�B�o#��f6�rt�e-��!�w�ZJe�����g�:��i��U��OiҙMY�r!� +7�n�NK�wBS���p���&�ƽ�YL���E��
���'��Qa�Cի��	�N/��'TG_*}.��u�RW(��G���{�6�N�_�X�H�'59PH.���t?;���i�6�p�_N�o��r�z ��R�s/n�#s���˾��-��J��&��׊k̃���( ���]��� aG6�3_έv�:�����>Zp��rZ�k��d� ���u�r/�e������(�9ٻ~����L�O���O�c�kֱ�E�f6r>Zq�Y��Y�H�AY��qg12ɋ���m?��_�Zr��Qҭ��3{�t�^g�o�l�Y	�Σ����JM����q��N���?����6�
':���%6���#�EO)�����;4��U1��5�:���O���_r���k~�={b/��m�Eʘ2���b�.U�^G���~��`��B't1��Hr(~�n���?T�����d)��M%��O� �Ik�](�(Ի�^�a���t����s�ʋ7��+�(i	��kU�5#6�~��s=`��oB����[t�8�*����f_���=�<f��2����T�%�r�?,s�"�IQ���� PR�i#��N��T��t�l��vO9�7�7���(x|��s�w�z!��԰1�7��9cם�/C�. ��:�k��Ԗ,8?�X��nŅ�F��q�� �*p}m����7Y;����� �Fr��f0V�ml"W���2 q���|������o��4������.Q�&J�e�.�m�kNo�i�=`JQ�P� �l��o9�P#葇]�`H���CD�B������Vkm�V��V�{h�����< HV�����G-80�i�v-,$ �^S�y031�|��	��=B����d������etZo/�"�9�)��㔓�/^��D�0s	ᰛ��*F�����~P2�x{���ɺ0rf"�4i����o�Ѻy�gW[�Ckƥ�f�l�jpgm��������g 	�ύχ(���;��d��|iۆ�����⩧L��s�n�ػ��>G��9��nS7���gH��+�g�� ��H�4j�HīD��`�[ɨ�� ��йY�I��9�W���#Y�P0�B�\���r�GB�.�3�ʥ_��4+�X��sl����
{덂�'55�WQr�v��/��!e^K��z昭:������A��~o�(��r�:q��vL��&4��[AԻ̠����}-��U��fD�����܍���4�FΕ�ձ*�å]N/f�H�7�Č�[�
F����������Qs8�p��X�%D�0�%�
>���dC�`�`�gzu��&a8Z�EeK-�e�`A���d�,���I�����~^E�P���6,V�k��U��9�-ޕ�����Ƭ�A��I��.O�}~�T��s`������ᬆ[+M�D��*�ٛ�����q� +9�_|n�������t�m�������<Q���I�	�ޛ�b��>����d���.�ݢ�xP����(�!X�xDr��t�;'��0M��a���y���{j0&G����ȸ��H2��G�������X��=�S?��E���.��P�t��?�56��s�g`��:2o�/RUH�~��`j?�R&b�<ڳm���xߗÃ9�����~������D���i���5�M� Z{C	+�,���<��:����WU�ɑ�u��PP5{�sQ�DTӁMZ9e����4U�{�iο�����E��ϑ���]N�b�A���[��B��B�6:���旣�����\ ���Zv(N(��o�HQ3�$�?v�V�6J�A�NR�f��J���oXs;��ɺ:6��Z�Wk�H�`M@�\��c�������4w.���Ē�K�Uvԟ��҉	��� Gv�-�\�T����$�+�8��nM�BRV	q1���ؾ`9�y��3���_�#|��(��/�7����)��֊9��p V��o�0jɵ����� L��r�|���I�yXg�>���<86��>��3��0tu�'�����A2]id��3�Ť���=h6H� ��/��<�WO�ײl2�ף��2e~+*o&�CP:Un� ��;�W8765Y�����y���u�u�HW���ݳk`�Bs�U����֣�Ql͵P�{zL7z2b�4-uͯs������[Pa�s�H��<�Y���~���{X�55ӧ�Uޟ�Ha �άX+��|I�^�v
cg���â��g��cd�d�f�,1tg�q�Z�"�)�J)��!�Q��Z���1�@(8�b��L�å-��b?��(i0���b69��dd)u�ҋ�|9m���]/&��m���l��~�6���P�����m�zb8�y�m�("���Y��,i� ҿQ,�/�!�%��J�m�$��L�����h�2`��Qf�a!�!�D��i�}���$8*���z��|��RJP�I�̆_������x~o���SĐF곴��!N�o�s�B�EQ��)�?�ilG�z���]�S�3��O�m��P�Z�S��y�?�슠��ЗE�$�q�8���e.��I����ܡv]n�>�u��Ø��s1���@�2v	8vQ�VWM'@C"�������C�`�X�Mpx��0 f����e�1N��lKg �00��~h���RAY��{/N}���Î[v$s!W"
��q)�ܦ��8¿�u"ŉ{V��7���T:]Z��.�fL9�����ۏ����-�z@�Ȝ��༨
*�7w�d�6.�嗩��s3�����]g��/3�l���
��%��Lѧ�̘��~F�'Kjh�R7�ܒX�CDx�x"}���Z�	Jړ|�x0aBxx������+��p_;�5o����6nH�^�<#�YǳrT�Hn|�op?)�c��g#(��ٵc�B�em�H:���0��Yõ�_U������-5p�EPۧ���1��h��G^���ֈ>�?j����� *H�� ��C�`���A׋�(H�,Ƌ���3�ڜ���V}V1�%�`?�3K� Y���r�����$��v��4�z�A�E�/��t��Y�L1��l�͞�m/��� � �=g�)�<�9�m}S-vf��f!G�(�D��u�����M���f�/�1u���	���/���2g;9�ͯ��uN�(�k�[��<�>�~���I�y��ۗw�V!�'q
*�X�G�i�FB=�b�Ց;� �+�zf���b�ԧ=��c��&bU��2j�4pDZ�e��� �%&*�Ƥ����s�:SJR�Ѱ9r��p3G}� ��W�����j�1�y�3��L���8v��H@*^��J*H:��+co�6��@��*w�`�U_8.c����W�ަ�YL�O2�Ѱ�;E�m�?,�C��!�e���6s1no�^s [f�g�c ��J�/����7Q�U�?<7���9��=&�j�> Z�6�Qe��;M^��*����m����5@�a�φu�Sy���	 ��b�qK��9Y���qu�}�au ]�7�a�y�چt���r$5�?*n,��]�̨� �*	���@'zF�0�̖⧋�Z<L��q��u��e_Hh�H^�ɝ7^ !R:�nx�w����эc|L<��<��L��u��W�sN�+�KmjY�GR��a_�w~� H��	ۏ����k��I4:��,���3�@�k]cG�7��U�j�t̀tq-�&�e�s�2���*.Ѽ3v��V*u��/��D��?�qK�\�Ϙ�}�_P0����A�����a�6�,�U�b��0ʕ��)���H��v!����o�;����V�	���a ���M� �<�l���2UI���Ը�P''_�G�6T)��WF4���s���Y�F8�1)緘��A�r��P��(7Z�T�ھ��ㄑ�|� ��ǧ����g��]Aǚ͑6�2l<)��3��8��=��<u�׽�ѸS��GH��� e)���I<��H�a��|ٖ��$,�)h�h묣<*�4I�oX>Ln	|,M`O��T
,%��o�|� �#_��*B����e�L�
S5���%�Ȱ%�W0��Z�l�+�p|2�Hک��M.���h\v`�}̱o\ya?#m��a��������ܮ�h,�Vqݪk'Ԗg��xڃp��n��T�LД{B�wnBϷ�<�]A����;ٗ�����zb��P�D�[��;����*�$!�Z�"�c�!d!_IC�P�S^z��.����90�b�O�jX�\�ƾ����@V[���� ���L9K�!�ꯒ���� w����rp���<-��7_ųc!?~�7�(������Fm�L'.vuֻ8��.n�����
�%J����Fj�?>�Q[�P$���Mk��^���GnA���� *�,��r���a�XA�2��ڊDϤ����~���z�<����e;b�l�%X���0�ի�I7��2T%ɰ��e�
'=��ۑG�8#{��<�����P�)D�A�Of��d�F�nY�:WU����������c@bE(aU7���a����V�b��*�u�ʬ�N<\p�]Uc����E��"e*���E�<�yv��T�c�>4��[/�ɣ�4�Aղ�i�h����|�\V'� �?�A�ݍ�/�����3�f4Z��o���R8%	.�k��0sy�8�Vk�$�(��x����l�#����}�L�U�:��ƞ�8�SYv�@�mXv$�l��@�Ŭ_��
M��Q����4��
��)�ty���ɴV��L����=����YR{J\�N@tq�6B����/�2Ӡy�d��8����>ʉݒ��9�� s�|+5��J���Af��M�����L�r�7E�s_ۻv�j:�r�&���wAw�ꖨ^'���ţy���`�vP�8���YW�\&3I���P�#t�0d���G���7��fÛf�2=n>�Ϲ��ǘ��
n�O�h�P4 �R�x�{%�]C�M����X`c��3�O��.��2�z�����ɀ��NسO_���lc]��l+;lYm��� �&����S���A��4���R�j��=�7�C��U8E7�x�e���LzX�F�",�k��>�{�|2�ݻl3;���/7
��X��Q27��e�	oxooҳ���/����{")9po5U��EZ+p=��WD�m7���ǖ��8�`���~���+ֳt'�S��~ղP�S�%P��q��P��Y�$>�=���R<�~-��	�:��R�r	���V�fF��$Ƿ����5[ZT��`D7��9s��I!�������uE�wָ7���N���G�Y�F�}{�&�ٍ�n�ٝ���DM]����r���X�H���N]^��#9�o�!D�LP��Mo�g��s�g�'�z��@���ټ���@�ა�G��#dwb�GX`�AV�h~@
ilȗ@c��?P1���g��X�g|	��ꁷix���avA%)hhx��"��V�
�>d������dU�����W�������In�Q������=����ݘ�'O� O���B_MwuBQQ�2EZsM����f�U�IB��3J�����sv�%W�B >ƋB���٢����d�2.�/�f��>V�&w�4��VCM)�P�đ�W��Q�L�wAۦk\N[6Yfm�F��{8O��޸C�Fy��n$�z�C�L�&TI~�y.���MV����ۛ۰����VT�����Bn�N�֕{Y����wC�r󠻆����:s�ke�?.��>�i�$�(��}%�5���߁C5���R�6����۷����w[['�g�c��ԞD��T�7�1?)���[���^��ȫ��NR��ߊw=�U6�e\���x����
'H�*���Z���4V��{X���
ՅY�vE����ڸ�8��Y�H���H���(C�lX�u���m��7��~�w�'�{�Ӧ��L��a�ȼ�x}�鯈���@��(:����M�@k�ԆP\��A!����k���Wg2:�;��i{��;<��f��Y�Ї��u�����)i|lW����Q�σC�og^��#�W 9�J�ܴ�m�����f;��T?-����*�,=ņ����WW�d�<��9Os��nJgaȑ���(�c��[��_�bP��5���!��.��R�{M�� u�I����f)�ft-�}Nh�>�T��9iU�/��w�-M{��j���&�Vgy�|N��G��M �@�(HW*�@!N�G�+��^2L
�zsM8�h�=�����G�
��ͩM X���J?�Xa�˱4��;g�菮���4�Ӵe�7r0��4��:��z�S�_�*^�=m�a;=�m�\�a�4eu.��΍�&��;Q׋7��/N���Z�i�X��>�X���}�c
�k02<��c��L�����dx�XR|z�$��EOZ�D��5ħ*D�8�t�x�6�
��P�o��ַ��S!��=״
�O��.a��Iʪ��Jx�dn)���e;��
��a���t�Ca�6
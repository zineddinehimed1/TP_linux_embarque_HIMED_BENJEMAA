��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���۳AW����{�u�)̥�d�pM�y7�w�1���'�"��+m����Ԇ�@?D.�#���A��ey^�??fi08H�w�%4|s�.���`cZ��wʸ�0�h!#k�a,�ˑ�lx���\�:f�2ƴw�Ͱ��7�� �[%̍�|,l:��>�O_� Aٴ�4ng��Y3:%h"$�h��T����U�\�a�,��@=Q{	�P,����=hBC�/�O��(�c�E�3]�Z��Zh�Y}�~���{pw|X�<OZd��Kb>�l���Iӹ�r���J۱3&s��:J��?��%B�G�I]�0��I��U��{�Dݯ�VEVE���Lk^�Z8`�p
H�#��؛�t}�lu�d�<�/�(�揍�ærY=��d#�X�yͶS�e�wXP�9�XG��og��V� }Ӹ^�����s��*N������_�e^چiq�T,�w�g}B����=z��Ҩ쪼�^�e�l1�r6t��G�����On�X�x�BJ?�_����/%�EO��6�lC��U�"7.�jrpN����`�I������t���k�$��$8 �g�} ��;�`�G��j,��B�}�V����5��K#z"�ء}��)7F�D�7;��*�m}(�Ṏ �氀�,�?h�t���In�v�|Ǆ���*H������Cf��B�B�p��N_:���H?�cQ�%��0D��]�:�;Dd!�s��Qh��m�Y�W��`@���Ƈd~���U�s�<�;��ӈ��B�RT���)�������.*Va����JM�p�%�p I;����h��[y����b��ѝ�V����.��^!����v�ʧo7�����C��rV��7H��=�qE9ar#5�g��Z8��L-�q/z�������}��_����zӥ���aDi��>�@9�h� BG.B
�جAP�a�Y�۰�d@Q��T�ѬnL��4�; �5ܹ�[��l��ʠm�ze�De]��.A�V���, p�Ŗ8=2A�Zvo��;?�l5��yq�)�G��њ�����B�&����䉥�ُT��4"-���P�C�t�L7՜N��,����"�mT�?�9]g\Q��.����JS=+���m�[�WF�",ڝd��ܸ�-�]�5~�����W��R1�@�`��6�z����_�|�+�	���R3��[������H�[}�����E�3ԋ�C����bz�>�jY9-@�dةj}��M�v)Ns�~Gn5�O�C	_��˟���%�iC����{��9���6� ����U�ñ9��v�(��Zհ_�2�5�گw��[����0��G��];�7�[�FB_��Փ+������#�J_ڍ�E���{�i�L���`�"�M'���/
�Y:ShgQ��0@8�Q��!Mh���R����wDK�����[*
w�c�#xU�����(�ʵ��*�в�p���y mZ;��*�HNL�����\�Šf�R2�����(�ot�pJ�V-�5���ߺ���{-�`��,tp���)��xbp�d �]�
z'o"��yS8r�vu��ň�³ߌ�2N��,����oE؋<@l
�c�<`�^�*���w��5{��+%�A����DT��ҷQo�2��ޛ��ws�0��Y��yA�*5����j�8�N�:���G�Y���|?��@�պG�R��ݠgՇ�$*bh3�����!|~��/�a�
T�)����Leۤ��>.W}]��o������o�̙fv�F��ᚧ:�e�q�2%���i�bL�vPM$�VH�n��]��_��R����vRS��
 z Yi�ZG3���a�1�'fq	�� '��	}}�����:QJH���7�8�T�Sd�78�����WH�p�[�w1!>���;{�jDen�Yv�j���a?te�H�ZH�UӴ�i��>�0�Ֆ�M�	E�H�ꒉ�-Zbދ���q$x"�}03�_%q�KWm���U�=fl�^�Yn����l<a�%��AnM�Q�1 �p
\s��_@u��	�j�6޸G�>)���)GS�� i��F���1�	�M����?���{�0n>2[��|L�MM�{a�����������m_��x;�k�oX]BA�)�2P�U�P�7� �q��Fnk�Ik�s#z�Ky��%��(>���yVG�6X���7萉���7����4�V���m2��i`�F���X���.�'D����!��|�:�����7ۃ���+-כN'e��v3 ��$���]Y�"/���S�;�4� -ؽ��^FSY��D����} ����i.q*��rw��a�k��<qH��'�@����bhd�(Q�۱6I��#�i*Ksh��Ȝ�f��H�:a�׌��k@yv��C6_�Z$��@G<���h9����^�-H#Q��Gf�U�x��/u�	P(7_!�aUi�x���~��ׅ��n6{H� �l��&�fCn#}g�M���d��t3_oUI����h"7R)*5&��r�������pp�r�(p^>��W�sv��s��{��a��F�f�M��Gi�q��_��:~E ��p��P���澛�K���+q�i��,+|D�8�|k�yl㕵�k�\�ȟb?Β�@]�W�����N1��M����i�;s��T��QO�M?>8�#�-	i)UL���̱c�#Y�`�r�Gܡ���kG�A��۬~۰�6��1�(L�xo9s���^���
F/ڞ�Rf�i�b���iG�wm{&��
ϕ*:�=:3�2r�Lvt�7/�B�C�'�Z��^�a,Zux�P7�H���jXM6Z^���zG��t]�a���ʪd@Z��j&��i��@Qʰ�?���K�b�Mo�������^^����>N[�,�fy�U�7F�C�;�]����:gb@�o��7$��v�	km[� �-���m��/ϼ�/�D�9�ϻ�u_���8dܫ�~��(�>{T��䈌��3h�?>���ؒ>��^<��~6p��>��4� �^�C I��D?e�V�� ҫ�p�����D���	&��s'&����(����F$9��8�0��s6N���4ݒ���اӅ�80�h Qb���/�h<��q�(�]��ɖ<�%��|�$1�R��b���8�q��������ω������;��uf궗�xY��m��`��.��TT����u����쁭&(��r�����{'��ꊡ�x�
U���{�V$ܽZw�q*�pT$~W��#�����aԔ!JA4�r�S�@%��;�
��M�/�f�U�c
���sVw5v�p��(�h����%���6�\�����a�@Q��_��!����͎Ϗ�:�i=ÆR����[+�`(����n���=�pI���V��>Y���1��Z���㊮��*�5f��c�,(p��X,Ӡ�v'�y�����Dn�y}&n?�d~��j�W��[jY�@�o@&���KHM��^�����J��b�T��|�ӑ����rh㲯��WB�R��'�:�|=��J���d6���Ҧ��ݶ�e���`�e=*�g�?ڣuG��q@�Ft����$T�gaclDuD��&�����j���F�Q��K�}���p���y�?���|Cю������-#w��?A�]_Ӥ��ָ����)�yR�a����/���n�ft�2� �pl��!Lb1x�"�BP�����q�5,�T���+���sl��,,���E �H��I�[�O�4�[>����4�k���_��bCi8d#�ʇ}(Q�vь�!|AG�1EN�<ѻ�I[i��[��~�9���QsS�lT֐T`�?yܧ���%;��!���=#
<%*���d�Z~2k�������k#��GL�ެB�b!oNo�#q��M������p[Aǆ1�Jw�?7j��QU3$�(5�;Nc����˶��N[Lo�߂���'�:�a<�ν����)8��x��(�ǽS�s1�{?��e�A�`��r�쪧���Fc�2�O�Rh�~:CL� �z�2��!�Q�1�Eۃ�<:I�����������!�P��5r*���y��B�g�4�>�m"���"�gɱ�u�Z�U���5sa�����0.z���H��V�F���׆�v ��$�)Í��ka�l"%Yh*Om5�X.�;1��C���^:c,`��Fk��О;���&:�$��U�Tې{��.�������^���丹��#�顧 ���>=�#:�	�X7�p0UG��}�WU����tO�t�d���Ӳe�� �X�����5[��l�v[��Pf5Û� I�s���2lw�Œ�
x��LN���o��6�}2Ŧ�9�$�7�� �w���-!�[��lW�86�[�(K��������Y;9�L�����p�!v�!�vC$o?�V�,�9Bw��4$��g�'(��p�7�m�}���[{�P�y���\���'�Lu�q2ѫ�6r���S;�+�E�V�il���ܣ���}i�����XJ�XA�����3ۼZ�G`>'��CaV����Q.�0$U;Y������Bu��Y�R׌;H�z�E
��[����܃f��e��BÉ�)�G�1���YW��Ew���Z���x}���9l�m�u>��dќ�.���g&z�4k]��0��S�g��������X�|=z�h6пHv�s϶[�7^�/9��-�X�(52Ĝ�$6��``ί��߆�LYqKr:>ԏE��V��!77����ᦻ��oma�~sm�dkXx��GJ�Ct�^/�}�X�������&���Q�c����t�F��I
���[��ä:96*�L&2����X�]ؔF�c���o��Ɨ�]�@?�ك�Um%��~
<��������}cr-$P�U[���� ��ؽW$G������)fl���B���U���<H���f`� ��b�>�B�s��U%�ǒE���s�Q+ۗp7��`���,�2 fˉ�eD�(w5�D�1�w d��F��ޒ��C��n'Zw�ا7�3���0Dd�����!���>)�I�y�P{���\�ެ��i8'�h3�>���%��;;{�3�����ZL��?�+e��b���Ş6Ď @j�`wG��=�j3��gM^ϥ��Dǻ�ޛR�#t�VJjg&7�0 H�~K���РMc�
V+ �kY*})�ww�#X�~�S�m�"x�@�2�)*c����Uŵ��}l��x��KF%�ѷkÜ�z�z����:�M3�ûV�J"�՟�^��c�چ%��ƣ�y_�Iا�:C��r�id����{=��)P<�rmA���關MLăt}A��:9��yƬ�a���o�"^3%j8�Y97D�k�G�ڝ��[ +Չ�k>J�ꖹ���ZA	�Y��l����e�Xo��f�R^%UNժ�=PFh*R>aAE
��hK������B����Ҥ}n�ZЇ� DE�6K�T��u&&����ߵ9#�e�"���)`%Ə�6����J(����羶
s����!�C��úŴ`�p�������ݪ�vU����+�69��EK~Si���B�����=j�7�����[�e$/�ok��g���
a��� ��&��L
0�e���u�M!J~d�
z��J�d���]3�9�E�*v�,g\`·�F�bm��ʳ�s�hZ�50��Ve������WKOpR�c(O]�B#<�/^���H6�b��o/?_�{~�|
m��:�c��P�&$�x�V�P F�"�a߇�$�$Q���#�8�����E7j��I?oub���h-(����h[ަgq�n�孅����E 0a77<G�F+�|�N�-�O�WZ��n�L�&��pȎ�E�ӑ��z�)�1�*BL;[���������R�>�4�4U�i�L�΁(�f��ߥ���KT�r@]�7'��J��v����/o��ڹ��pZ�q���ƓQk�3TI&b��#��VvyG>��y�'k{c8�Ѻ���\7d��������V��p��oQ��3�F�Y�X�2y�p�s@���h&���5�^��2��XON�
�d�d�r��2��7g쳂�\��}2eS��nY�t������ݔ9'�*7HM��u��7ؕ;����qmQ�;x ��e\�Hs�ڢ�	(Dr~�]��3LS+��\�z�I�HY(sk���	�M&�	��D����n��b�|Kʩ
��z��?	t�Jy\I�C=O��t&���o��Vغdl������/=�}ӮQ}�4r��&b���6��_u��WBMW���Z�ޞ`�r��Ҧ���&sA�z�n�M%�Oof�,��J���i·�T�5��Q9|_�ND+�(�N��ZR�ZNQ��A��x9���`���kO�g�0f����[�-?B�,t�:D��8�C,�<A1g�ݴ��v����Q3�3;��w���꿄�_%���g�țHR��;ۧ��	�i�G���6��k�i�$(�N�U)��E^�aEOf��#�!q�}q8~�F�>J|�e釺q8DI���.٘g�r�o� :Q
�vq�����ڹN��*n�e�Ns.h�{��'儧�I��4����P{�LN�MfI+V;>�Er6�ˋ#�a�U�	���$�QC����Ĉsd��Kk�m���Z��!��q�4���ZL��k��z_q�@x���T�%w�B�j�S-hv8Ih�_��Y�!��"QPw᷶���b,ا�Ò�d֜�-�s�Τ/d���}�"F�Ty�m�>M}��<�m�q���J�:�$6���*R8U�?r�������ďd.?�eO`vw��z�V��x*7 GW� �
���ynE�ʳݸ4�L�/��o��4ڮ|Y����>�[�ǶJ�z�VC��/�7�%��k�2���}�BCW3��3�P(��n�5U�"��+�q�mG�	�-Ԗ6�Y��Z��LϪ"D�!^zU��ꁟu.��Q{Q��`J�� �|l�U�
���U��`�wq]����^&*��@Ёﴻ�R�*�IDs���1ʬN� %CS��U�FZL�������g����:�a��yv> �ܿj1V�<@=9�c ��Ե!�Bo��6��HJ��36��ѓm�j��Z�F��� +�����yJ^��#3!��'^�;�
���ĵ�2�o�d��z�0�聞�L��x`6l|���44�G��2��n�w�Y,��C1�lN�P�5Eؖ%z��Ҧ,E/β]L��k-��ں���uƏ�jp֦#E�H �[�f^~AY_��q���Bcd'�1� g>�\�ƀuf�:k����@Ee�޼%�X������:]�f��J �+�1d-�0���Z��Ĥ��$ݢ�|�VE@�oI��hDy�
��`��%39uFKx���|6���#�� ��[�ŵn����j8(�� �禅�C��d@$���Y��E���&�:s����r^���Up/^����W��D<�n����ƾ����2d�$���FQ8��ϸ�������w�^3�:�����|7��]+����l�h�u�Mj�R}��s����g>���~��J����wX���}5~#9~��t*��I���5��o'>ONts\�|Ʃ�b���H��έM����t��Tǌ���G
.�G�]U�9ћn'�1�U�߸�[������U%� �����C�0�d(w������*6�8��5l�L|wU
�叉cHz�$FJ�I�Do�?���Į�aK>_ῗ(�9J����*�)��Xc�f��Gc��R�H��.p�!��:�匄݂��h�m��.��U Z@'���F�#�|H�	Ʉn;Vr��<��	&Plǂ�j7T��P�t�<���D��i��WOl9`�M�=C-Xt�=�nV����|K�v�-�]�<Îr���,O�3=�*-�U���`?q��;����I�9�d���Gv���@�P��:�)LT��ԟ ��3�$\	���:v�T��
�l����/�+�EJ�2�Q��&�}|�D���V��]?��:���zM��f�3�7���J} a]nB�q���?�m>*���M��ii���X2���~t��}�7�M�U���)���4	=���L����h��5i�t��W>T���~��Ds:������.(��AF�w�zy�ǐ�ܾB������x ��+7\F��I�W�nY� J�L�֗U�f��T��S��"�J
�߆��ζ��`�b�9�^m�*�
�:b3���6��c> �C��'O�x�(��N��?���$y$޻;c�ܾ�?�V����u[��ⲩA+�d�󓙇�B ����A��g�<�+�6����;�谍�:��1q��r�����,޼oZK����4I��v8f��$�6���H��{q�v���f�ߧw�����K�I�y�|g���18L���W�!���d.��ѷ$0���D��d�S���t� f����ׇ�I@�!�n�uՃ�@c��ę��k�Z���	���Nʄ�Gw':��p2+���	���o$��^mw3l�,����ꆳ$��{�����DF��%@�E	�!c��E2�8��A�Oa�m��	�M���`&J3�����ۋ���ՠ�/���Ei1 ܹ��&WJ�k�Fqf	=0y
d�|���U,����sx�J���V4��Y\�>��g����4���#ad����B�ϯN�ps\�S���3�!	y����
��Z0�M@�2��Ja�,�����w��ͅVNx�3����4Ҵޡ&m�n?���0���ɇS$�F��P��e Z�ߍ{ر~��z�|;`N�O�\ZT�e�����xxZ�Y�5F�L�i:�0�����j�(v/!։#�W�-ȴfw^ݷ�u�7�.���Z�蒽�n��D>�W �"����4r�%ϳ�2�����������I�,�o�%/ E�9�kE�m�;I(K�_u�'.�"�H�~��z����4$��5$`�����,�%��f���X�hCc�=jƩݞ� .��l�Z �vM���K���i��e1��z9���d�(u@������:��.a�6`[� �c�8�_ߙP���T�6]���b_�~�.C'������m6^�t��V���<,�^G!��<�!�*f=?'���_���9� �v`GL� �Wo�Y��u�w��e�Y�,x\���.�q�c@�a)^9��E�Y�֤kH�?���*90����/c�[�l���فJ�?�����������Vz�d4Ae�SwwT�A��ћWT��'��MA��9�VqL���e#�gT���>�{X� FJ�2�|�l;5ɞ7�j�H��8/3^�݆Jֺ}eo{�fA͵�bat@xV;e���¶��r��}��W!�Bd`�)��;�(��F��֨ �S�c^oAycU���c�����ϓUq��q�uP��P�|�R�mw�g �FhF����^���6b��ɠJT�n��#T��h^�F����NB� d'��A����?�[l�_{$�������Y�!q�I��y`>�vW%��'�~N�L �>��`�EY�o����mЫg���@z�{��ɾ�VഅKi�cU���>���G+�sד���[�o5lP��L]����\DUǕr�˝�W�@~���^�Ul��������Oa�]��ƢM;@|-+�J�r����� 0����nje`���k�8qjlK~�:�s��>����Y�ʫ3�PӜ�g���9����l�u�ʙ�tV��`�P��Af�xh��F����զ�ѽ'�&��$%�n��N���QZH�+t��������7S.a.џ��np��F�c�,g�`�����C0R�s�u��c{D�����ɻ��/
K�'9hc5�a`S�Bly�^�s��F�mJ��'>�5:�s��� �J�r��>�w<�E}٢H	Ut���\)�{`\�ᔿgQ�w��V;v���q����vEs�Q�0r9�bw�3��'�k�����M�a�!�� �{L�.�������'��\&0�S��H�Gw!ň�D���N^*�٪�v՝6;T�K�^�Xv�í�M/F�����˾��W�P�~	]�[C�o��ME����u4�V�Ec4$�&D��5pt�e�w����z�uR�:���Nn�U/�Θ��~l�y<�W�%�G�1����;K���V���'e�� ����o�ᓜ�\e]���xQ,���f���cd�v9˄U���������[(�'{=�YJ�s�9ɢ+�Uם�����<;��gЕ#8K~v��l��cW��n�찭��d�4ۚ���?��)����������cA�n)��xͮ;��όQ�e�l�.֒��N5���L��MH��W��ޙ�z���H�e|*�h�#�l���Go#��z�,ǕN�d{��Wn��.�rP�u�`y�^K�H}��[rz[id+����~;��e
����	r'+o����OHHb7��
Gb�@Ϋ��w	��M]����h���osD�]���v���yO�i=}+�}��n�f�hh��w?U0������FiNV��x=��^A �Q%ў� �&yw]��&���.B��i����%_����nF��X��!q�
^����qp�2�rW�;�bzz�J[א�T����_���'��?S�q�
	W7���*�18~�.�ϟ��N��	@�^���� ����f�Q�^fάG���4�R���3�5�����7�6"��|�������G��,�0L���vW��ѵ�����^���(?(���	�N̐/s����A���-�*1k� �(HR�G�@�,�I�2��Y���$L�A�$+6��^W�*���ƣ�)ێ T�~�_��OPsԚ)��Bb��m����Y�k�S6����!/P �i�s'T��M����Lt)d����*��酉�Ћ��e�a(�缸:5y���](��۶37�i���b���]ӈ�q�� 8��J����q����1�,��OeK���\sL+����XF��z��,�)A�"�s5�;���vr!e1��J�؟�Y��P�@T�z6�4���*\4]�ޱ�=V%lb�ŋN�u&`�ddT�3�iB�q�����i�V3r�
d����#�ߛ�'aWg�O|�4��zYq��l��L�/��='�ӟ���9�k� 7��A\���;�F��=�S�B`�B��BL��B�ˍ���q�'Cr��C�®��F"�����{�x��c��d|�����!���K����d�<�uA�A���������Q�fSQ�
�2/7<��$�Z�8����B�G�@}!� ��9=�S�i(
���DK41,���vYy[sm���������/́6;�m	���c�:����:��Nq���{�"�i�Lv-�ʗ����lS�A�R~x�jVȎ���f� '�n�����ce��,ZT��1��� <�x��t�I7���=`H�<��Oa���T�YZgjK���h5o�No�{����rZj��ϛ ���Z"¤}e q(�h=JD����ً���m
-xS�`�H5�,�J��پ��ߢ2<����Ї�������uo\��cDS���U%5� 2R�I��с| z9���lY�p��6ⶖ���3����������!�g���F��5�_��K�Ys�{�,gS�����KbWp'�!���`Er��)\��߯�75���"\Gt�Ѕ2MwK�������������З?��k�����������zt;%��[�5�Sr��v/��_\d��`�L�m<��{��fƶ�C�8�Pt�Q�)])�#��I4;d��a2�;`��� 4�d6� �,�8�;���
��#]m��Y�P!$p~R\����;�
��NA��L�z�F�ee&n�܃8*�4q�M�~��{������J}�g�k����	��G���"IƷe��ͩ ��	F/ڔeB�p�g�*��]KS���ъ��Ee��XR��\[0����ԥ9.�뷱�AB�Ӿ�w]:���1��'=�t�N����Mٱ�R!��>�\��������8�aG�2�h|��aK�"�H��}���L[�UG�2�Ck)� �C�4
�%����O�vl*_WVvozfY���9*������#)�V�Q��*��9�xn=��*N7�� tڢ�` P�ʆtɡ��D��:0Di%��k8R~O
I=��@'�.S@� �^�ӡ}k�Z� �����%�S�60# �ã�L��xw�
	�hU����Q
&6��������ol��(�	ֽɑ���2�Q�@�ӱ�������F0�����b} �rN�w��9x8���jdD���0*5kn��`X��6�[7��];T�����U��p��|�ߡ����a=��L�d�|��nL��#n������!f	�s��+��"��}Xz~�Ǿfzq��a�p1=���\�y���?��85AAF��DL��(�5d3�429�6߁��	����I �jSQT����]��94��G��Y���%I�W��w36��dѼd�^׮=�Fv��P�X��#vKcb�,{�Y�U�� ��M�����HL�)-�F��^ӄ�񱹄WmMB��\�s�F.��쇰�llU�0�r���ec��Ƴv���<���wfR�ss5u}n2�5N��b���g(5,�B�i�
�<ǥm��'����G��Y�pKf����;Ø�ɬ:D���g�Ȧ(���>{�ŭy7Q���ڦkഗ�S}���sf� &@T�m�k[��iĶ���O��"bg��	�t�y�೰��fV�����: z����@v��쿲�L�����v'o�gHLe�|���c�X�ֽvlf*�䳨lO}���'��Í{�}:[S�
��C�O�j�ǌ�+1��p7l��;Y�5A�o���s7�Jԃ�C��}k��{C�ʙY-q+���|l�Gk�Td'��L$����K�IrN���$w�Jou8~ ��]"�|�O���ΰ}�>� 6����������z}��9Db~ML�lV��M��Hq3��!�ZF&$��F�_@��]��Q���>�H)Oc���]`�}YyaҼ�[��Z >�z���i��Z\�?��|#��m�d�L�S� ŀ��f�7���\�m���h�aB�x+2����ٻ]����~��w���Io��<�si��BK��j�
A>f��2*�RKG5���xQO���7:�'�������w��#&ဃw�e��dIi��ڈp'�����ODf&�b�ͱ4�4i,�Sq�B���Q�����L�h��52Q#��'x=a�����5�v�i�DR���ޞhӱM!��U�F�s�X��n���-" ��1f���5Erx�? ��a*�N[q��(��WY)����Ƭ��E�9O����d�zKɑ�����۠Ӫ鍂�0z܄4V�����լ�{ �.�T��l���\�
3BbQ$��ZW'<���$�l�T�Tb�����F�#�1��z�:�b)�9Wx�ױ�8��I|3=w��s���=����!����u��/w��]�9�XB�Y[�D����B��WV=�o;�3	x87V�H�L *�l(?�.G�M������@�#J�^���Q���5������H섉���&'}K����M
U;�X�!9����}�l]��iv+	L=\��R;����zרDԕa�=*�-~��K/i�+�(_�R#�����	=���{��q���8`y���pY����teTO�A%������|�����n3g�⇎�2���qK<M�h2'Z�	�-���M�F�m��1�@�����M=��K|}E�J��ч0�s��hbX?\��B�`eSZ,�m!خޯdTV���+u�Go8N?���rWh\* �u���R����oR!�����E�5��`�_m�KSc%qF��8p��`Py�u}eںf�D�t>�����9�pE�����ل�?����-��v�&� `��b��Z|{ �@>��H�'��,P��n��(���WR�ѱg���X���R&7q��&�������vuJ��j�����;��=���BM���rIa��͌��P<�|۲1���qH�G�G]S�����r�m-ͽ�e��I��� �⫫ߺ��(�{��TRu�=���*�km���*�cRo�Cإ9;�~�#�_1��,@��&��>
$R��ڴ:xlP�i*9��i1$@D��/tԇ��
�1��쳕-�h�̿ssZ����2�*��+N^(�=��\��x���7��mr��żDL�B�����|(&]��Tu���Q1��H8
\��|wZo��c����SG9�d���������ަ�3M��^] � чt)y1��PSЖni8"���VY�(��X�Jrڻ��c1�`��x%8v3�ˎglRX�,�㩦`�x1!���u_R�_<cU��3'Q�]%������.�'���T^ft��ŊHo�2:�v��0�
]
ȂP�	�o�.�y�>h��ǱP��+$���J�����}r-�^A�.N#`뽤� m�����b:���I\�]6BU[��1��"+ �Q/�r>-���[�����_������M�@8��0D�ҁ�Z.мv&��:�s��zš�x�*���z�K��^1���ve�;v�Tj�D�ivjxgg�)�J��	����،g:9_dj����[)ٵ�_��\��r�Uܤ#L��F�`����M-ϼ;�ɴ������|�j��(=G��p�&�Itp�����=2���9��Ń�{|��y�!���r�n��nΝ�L߀�ma�k���uq�-"������������Tx�6�	㞰R���h�"q�z��ـ��ڷ��X�<�f�r�S@	�uƿ�8��9\w�^��z��1�;��
�]A�����u��a��K">.�����t���pX��	-ժ����dX���˲����ܩ��&���B��V�q���{�}��l�!���&0Ӏ��X޸ �K�tʈ�А���?gb���oP�Jۭ$F*<��}c�x����l�y�������a�GN��t�Df�:	\��٠1:!���/���d�I�Ӆ:�m���dK���8�F"V���7H�5Sgi�#�I�Ϣ��n������^�-O��o�/�"�n���
Fa���V@��E7�Ru�� 1��<������_(�淥ebZ�h�=W� �_a$�X��]er��`�;�vɇ��h:w�d2ɉC����
SJA�[��B@�n4S�
�s�0Y(��^5�gk�.8�6f,���Lr��!�o9��0�d��!��{>���L��h�"�~��ړ��-��xr]��C�~8�F[\�� ���1����o�%b�
��t��`��S�p�Ȁt� ��)5l��*-+��p�X^B+F��-D�!�|�	G�2���s
D���	�|�����%��W醍B�Yb�-J7�����zf�Q��(<��G���ko��U~2ޟa���/��'5s\\���"��Y����#�<���n�\>����jk�o{3�a����5J�:��������Ȗ�=L)��L����^ ��M$����"��ʩR3K���{�Ӊ���h:۸!�����)�_#�Op�n��[�p,���C|�<��`��$�:-ڭ�C\�8�g�B�hK��#[� ^�7�P��Ԑ_4�<�� t�G.hw`z�tL���UJd��>E�A���ə�>&�ɵ������8q�2G�"�4G����P8*���_, qg���`�M���+��=��'S��p��.�f/σ�s-������7��i�i~ŮA�1���cF� ez�#H�7'��M7{���Q-eRQ'Oa���()�c�uA��:�߼e���0ܓy�=0�:���og��]oZ���w���waPg�gqG�|\L�����TT����D��
���X�y��P���]����h6�V�����V`'+���Vt�Y_�]�0d���(x����F>�Yo�}|����T��d�o*�i�yk%Z��t��9�o� B�Y�`�z����n���A^W���G�\g������g2a*��$8q�5T�U�����݃����^	;�!l���φ9�u�Hg��/�N��-��4<-��Z�W��W;��u��;>/��K��	�U6z*���[i�[[����}���
7�Ka[����+���O����U�.J�ǋ�)�֌=�e�$�r����2:\	$���vy9���=8zTɇ��MCj�y���r�'��z���[��g���K� ���"�*9�7���(�A�M%�O�vJk:J]±1�m���z�(��`�/�syyj�ϸ�d��,�!z�ajta������ i�� ~¿��VA�D�>W�R%l9_���cpru�c�v�*MrG��˼�l���ugR� F���gP��;��N�d+���Db��6YbV&��D��)�Nc�eZBd�~���i,����۬�F��I_$���]���`Q���i[�fO`x��n�=6B����c��a��T��6�F��o5?p2ѷ�)��'AF��L[�;V�cQ&Y���1�]����DD��V"B����7z)b�|���y��|dhw[�Xuo��۞�h[/ i����=�ҡ�!������Z���0�%v���	C?9y[l f��\Q�0n�PΎ�s�P�D�$w�n��܁��#��5��]�d�z%B˓��y�=&!xv7^����T����^����UC�8Z	�/��p��R�����Ua�0q���@;����줥S�R�'��t̯b%���)1�O���n�Ǚ���qT�z��+��F����y��!٣�r�8Ŋ~�ų���N������������|=-�e�Q�XJ|B����WTL{� �sqc���v,"�r�wP�^��b�y=:3Z���:���xP�oaF�aLh�PKQ���[T@���/nT&�<��u V��0���\q��(����6�3E�ɪ�˪sc0�}v^��O��;�����*W���9lݟ��2�w_��\�&0��S���G�Y'�"��bZk��(1?L���[@J��%ύ�r�ѰV��&g��G�,=a�&;;����[]�DM�#��tm�I!-�����B$�EW��y���&={���+ƕt���`�t��d�O�$��M̶��iR�U�B~$!����Ѧ�����#�+�UD#o���3Ԋ���C�G ��wov�a`������8�p	�A�C���G6$����3���"�8µ	p�Iﺀ�)��/?���,!FL.�gxiT�aąF����A�����`� ��]��0�[�@~�g�m�w;FU��"�]u_Ł+����#�����`�?0�LX���𼤎fy��	��X]�)�J8ʬ�Fm6U\���j��ِ���(��-�7��)��H����o�Q�ؙm�S$����,����/.�Z�*�z��_��+�d8�3�|S��Ï����h;�uKKb��s.~c$�k�Qv ���C��T��D{��ސ�.��B
�i5.�w�T�ñ�&��d��|D^���0�Xw�
kjݿ�؜�Q���ǒ$�P6D���k1�N������t4ft�"�Ɣ���A�,������'{�IN��S�b�	 ��^���}���a����M�l"���k{ǅ�s�����o��bE������J����AY[�G�����@s�:���#
YO/p3_�%��G]9̶�T���D_��1�tV.�A��Y�������$�ã���X����Y��(�?�v24�'�y��\�o�s4��Q�c�?͔G]�vhH�4��2vKUyz-��N#��A���D���ra9BIe�t��+�Q$���$�˽+�	�S[�r��'����V��.�?_t)�,��]W�;$=Y���n������K�W�K;_lIK�N�b�pB��X]e\"�/D͋�?tS��AV�tdYΰZfQ��YI�k���o���6�z�:m�K_�L�<����35J���:������ tM
Z�@<TQ���{ �$���#��Ygx�Ƚz�^��9����-� ��Ƅ䯞 �-����{�)��Р�����w[X�*גQ��1� W�{��#���p�3DH
!�gI6��H�m�a��p���K�S��LtIF@ܽ�4_��c���M�O{��+�Z�)�Os����Ĝ<���w��
��E�u�B��Q� �o�r�t�5Y9����-�22%PF���*���@��*RL0-��������[��� s~͒ū�B�b�{I�0Z4p.���6Ǩ�xr�K���D�AףUO�fC(��]�2��  ��A�=,U��k����f�J<�}�r����#(����R),+�93f�&��n����G����q�p,��^���m̪Ҍ�gѻ�{c#���T���%��Om+R��ǝ$�+��f`d��gU7P�dӹ��
��A%�6>�n�B!Aٻ���Zb
خ}�}P��y�cL���#������=�kQy�)9-��Ksa�zl5�m��z��|۠��* �n�Pw���}���5{������I9��0�,G��MM76�!"hD2�D����O�id�轴�������l��;q֢op7�ֺ���K��Nf�$��Z����C�k�A��*�����{M���N`c�����53�f	��g��{{�%ڭ�Ǟ���U���L�=�>��:�b��N���Ȼ�7'�F���������6�q�'N��۪����<���4e@hA���*d��y��d*���Ю��K[��R룳h�s����NS,V�}����O:7��w1C�~��Y XtV�{r������}��eSw(Pr#��%�-�4�[:FeL��H�/;�k��L0�2N���b�)�$�bG/���z*rn��*6��YDʢt�dG��d�v|0<.?,����1l,����k:�7-9	
���^��{x��$�<�L��i/4�����g-7�������Ԣ��p���}{���[IO��u��C�M����$!GQ�K�.b[�N��~�]�����JT�{0��.�_����̊��+��[�H�⮼@c�����I���h�k����/��-�;����̥�o�fA�{R�},=:�P˞HR�ޥ�Q�%�h�瑭ߦ] ƖF�&nX�]�1D�����_u��/u�[��֗�������7[��|�b��*����u{4�g!*s&dY�R�/Um��񟪮� V�ygZ�+SBcS&bkUV��a:�}��ùſ���%uU��F�3��J �:�cS���j(*�	�Iq���#�5ֵ�D���T���IX�>�F�J��~
y� ��哄�f��z�XA\@#y���U�Pt�z�_�-WO{�z1��I��4I�sJ�򵀈�)���!L,	6ͤ�[*�Z�s����OPQ~;�2JQ����XW��C@�s�S B�$r��#���!-��/O��NQ���f�Q=�b:ָ�t$̖Բ� Rգu��D7\���'�9�Mޒ@xe�)�_ڕ��1$��I���?EwGh���uW��`+�bC��ɜ_*y7�,�;����~8�b���*���l�BF����aTx������ۗ�:�eH�����%�Z�c��-��������F%SL�b�U�B�Nw���0 ���(��1kM��z!�Ƈg�ɠXy�Z������� ��H��&A�:��e1��$d�nzVQ���؈`k��۔�"1</=
S��4�'�Q!�\f�-�

�����Q>#]��Pt b�=	F�_ZhEI*W23*sy�.�9V���q �S��ylP��A�i�#ՙı���@�)�,g35�:�|��\�L�?8�B:|ju�Y���٨3�]]������SΌr\�%������Y�9%�`zN�Y�f�sE�m�8��f��J���N�y��e��!�#��%��Y���\S�r� �0��\L(�Ri�˴���G�##J@�<��{��Ȫ��\~#p!Z�i���_��{���r���l�,��5`��z%9SVx�6�������l����@�'��kTL�ͩ�7b�}pzDz�0������Px,�tF�pG��U� }Hk��E�U��� s@��fܨa;�[����g�~4& ���ZLi��o.&}y�>N{�J\,Լ,��ä�}�W����Ȓ��LW�gr��I6�1ф�	t)7=9���4
.�<h����a��IY\1 ����G������@/����c��$���6'�e�A��"�;�A*��wW;�l�~A��4�ņEB,��4���41���t����sub&�O�4D�7�y�+lۅ��^^2�AP�1��UPE��ǥ_8*��i��.���Sj�ؤ�Ø���b�Ȑ��o7qҮ?x� +辫`�̲P��C�pl��^U�@������-Ŭ�$8N"]x�7����#�W0��!���	썺�7��x���D�!Hz��B��Z>)�\������M>n :�-�� ԏ�ʞj�������=�O�I��޿�:Ǵ�"�`�\_�������Xg)w^��^��D�-��ec����`h�<ӕ�&7E�F�7���i�7����T����G'q��?\�]Vt?� �?�[-�w����KW$�ц*�Ջ6vV�!� �y�Q��oL4)��#�y�*����Z����9аQ&b�x|�l����Q&��	��c5�S aa=G���{e�S����N�L�QI;@��=�	$���O	������Z��;V���ST�Ȣ9�
��)I��v�W�z 9�2b1�i�7�2:Ԛ[l5��"�܊
 vZFm�ż"��{�l#n>��^�^����ܿ�n|�T�|������Ao�P�����NM��̨�J���E��R�Zu��Ep~c@쯢�W�&nȹR���gZ8]�:U�iU$�ƨ�)`s_E�]�?���BТZuT^W�h�6)+K?P������l�!��P��3o��J�ڷf���LٚXUnq����a�\A�խqV�4�L�r�����E�@�qR��{�B�晄t�"H��}K0w�"�W0�'W�E��1���J�M·����C��z"��a�����-T-#������|r�'��-��5�n%_EK����3\����(�`�.��A\�ٮ�o��=��C�(��k��܂����@x�/$���D�ɕu}(5Ю�-�(�X�{���Z���/�/���el����_�&��r�|�*t�i&B{������WE
a��<`ȭH(�Y[>��tSsU�/b@ \��1F����t��ᰡJ!���;�ρ�gV~��gpcp.Rȏ�I�P?Zݬ����E°�:~���>A�R˿�I��1.'�����]b��"�_��Ū�����"���v���'Z���%y�k �wt���Xx�I?��i�S8s�2n"����Kv�f���}ߎ�;��7S5�q�SR�QX��&���6J�o7���'�>ڛ��?�J��,^�SU@�jN`}ne�1��6A���+��`����;��~V`�̌1� !��F�&��<��7��W؛��������8�E}��ˈfkҿvZk#盔x{�TO��v��Zo?4G�B�8rf�X�V��uU��	���JWTe��:D23�|4N�����>~��g
[��4L�G�~
w���x8%�O ��v)Ul��В�\A����jJ�65�K�R�/Z4���� ��0���P��J�1��>$5��[!�u���|C*4q\�H��@�&�R��|�����f'��@@��-��`��}ܰ�#���������nY$���HE%��^{����zח�����P�n���嶙���U�@�Q	`��ߠJ_�t2�����I���᧣����Ĕ�H	@<i���5Y%�ħ��]I��6�p��
s>�WA*�z����{����s�~����l!1�FI� v��]�-�ox��nh�bP10G��<����|��x����^t<E�@~ZA'ϒJ��D)������٨�G�)J�� w�N�h�l��&�
���2����1��gI��;�l�?bX
���?Jŀ��_C\p���E�U�FklI��[�-\�M:;5��L�j��� �Uh�!�bW�Ѿ�����Ml�O��=��\oCt~�i���|H���|�|Ș�ٞ��v�	Sa���q:��X|:Ɖ	�������שY�Q�Ě� �]² �����#�q��53�B�O�$� �IfJ�f�w���I1q#� ��7f|�ݙ�$� ~}�%f�ٗ���*H���EHf`��a�q�hEŤ�|n�b�a����367(�*�@���qY��s�
R�MY�&^.+nTĈn$s�([k#>3�� H`T��?F��sQ4-79�d��M˲eB����X���N6�6?�6��˟�i��
����3�Y7�~\�O�F:
��������H<�÷�h�B
6Ɏ[�����88�r<OQ�26	�f&B�n^��� �S�L�R]1��G��R9X�Gs�%�^<�JKISS4O�0*r��f:��'�Z�D!�'PЎ'�@Ί��?��V��D��A �W�����I���I3�!�%}�O\���r�&湓VMezS�̰ PZ�鬒M�~�lȑ�<Q6k�!�[v�}+�T���$�)-e�7��HݡĻ\=}�L� �A����e�����V��.�mS X� >>��̧�9W���3�BS�8�[�NJ�NC<�W�����o�?��� 1]+���gľn���=�%Ɋ|ytX,��]���p"v�'���|1KfSDȾ�Y������4��$��$�r�'��J��B��N����i�|�2RxSxj҂o_�4Q�ɐ����	�R_j���M[�)�u��+�D�r�Kn4Gd��"7F^L^�@b���1�0$r��i�(N�A$c|�d�x��k�z���Q�d�]yJ�$C�Z4q/�����Pa�j�A��Q��CB�|�ȅ�QZQ��Ip���Ļd����="h2��ucQ=a��8����0殺���1]?+�A.zO�/�<�g���,o.�>�5�('�������t����1y7j	s���e�?"Ϻ�����6�2�f�}y���Ah�i��Y�7�S5��N�M�zl<N�+?n|�LF�|RV+��)�ؿ��b*�1�ϻ��i@�9VI�5�����,:ׅH��{8�X�P[�6r���?���[EuC��a��ϑ+���>$m r�PX�}.T��5i�=G�_�+����lN ���X0B!�0��u�k&�O�Q$ K�ke��X�Ѫ�V�>�G2��G���' x��LZ�h �n�o��Q��d��l4 �#s��w>�]�9 �z���@����AY��܏��ƩG/�V��5Z�+�4�pƛ�r&x�0,j��TDЉ�p�5�r���gh�&�9�`�;���t�h_���;����yT��.9��z�\+<(;���F��3xa�KZ�k��c����Rjp��NR�5�7P���7��L�stc3���HK-�����!a	�:���FQL�l����X��f<�o���\����ҊS���c��bs(�8�+BH�y�~�6A /E��'�o ���l��.f����B�2���5+RѨ�&�a��K^s�*��Y�4��|*����N������o��R�t�g4euS�	���.Z���p/%�fZ���Mԍ%���������b J���R:��1^/��0���^��6��bҜ��J+��.��b~t"�rO�#ZJ�B�RQ��)v�1/�?�fv���]���K�a��nc0�gD�طVk�A�����!�15�Qb��5g��Np7G���^'���E����f��2\����W���dpg|����y�O��1��r�w��b��T׫Ao�A��|�?�d+6���k���ʮ8��<n�<��oǏD����S[�}�����ش��<��\�D��x�r���BR�3(�(7E4���K���[�&����d)�E�����5��@�1<)V�mj]�]��gBW����!�������~�&avN��#��X�\�}��H�~Q0�8�����䁡��&���/�^ht�𖒬�dQ��ŷ��\�O<Em���>�NKGzz� ���#&0B���\w՛��J��A;����	$�*N��]�g�Q�B)��=&A$&F*���AY�T\/�0����y#VG�J��y8����	�#��vY@.�΋N'�3-��S�6CBs���$�)T��&��j@T�.�P�>��8����lGM11<�m�q��	�����u�a�(Ffc�_�cv�e%�&T����O^��$6�)��Eo�M���T�goE��R�v��☠��;P��B&S3�l(M��wtlKĢ��HT4�������~�)�<1"����U�.�djB͒��F�*tk���qj�D���.�H:���0-�N�q�������M���	O��e �K�zb�!(��-��o�����H��[��5�V��*�
���s�	
re���V2}άs
,?��&5fY��e�f�Yʋ�PՖ 
�K��!�a�t�pzP�A�<X��iDLA�}�&��m��^H�>d����^�6R����{6����*>����4G@or���o�x�]B�������%���kNJ��&A�C��o�"vA++^�3���;Ov��JlN����?�Ւ	�w?����I�~��qe��&zeV4s�0]4� �0��7}Gƻ�c��������d��f'b�_�3��Z��#)d���� �q���x�pI+������CyBv��+������'��ϸU��V�� ym�)�>�
N�$���#�s�����D}�IU�Nyx�'cZmГYY�
\���(�í��w0��R�ò��}�=��
�$��<6joI\��?��K�2}|^�b!�fe��6gM��0� P��� �!ƽ���p�YYAJ���*wa�߮i/Ӽ�7a��1G�т�>��z���BE7�\�c���r��s�"�-��n��8��'�T�My��=)�'��$�̀�3�9,^�Lq 4����RѤgH�DÑ����e0����#��y��@x�v��M7�p�qYyM��(Uɔ8<�U�F����Ơ�q��@F�� dvٓ+J&n�97�-����J�f�e������:���-X$�(�-�,��g�(��@D�2���!�
'7d.=\$rq�6� �1��v�`aGگ��~����������3JIYy��M��l���e�Zt2�T�6��;*�(0l�oH�Tɥve�>>Tm*�?xk�����M�4��M���8�_7i�oߋ>�|ȇ/*寷��T���9�=51��,���4Q�,gK��{���ʀ�#��|P'ME?ř����Q�3��#���B�01 ��A�oW���y�DXk�������C�F���7,��p���8h����:팵oC����ݴ�s�I}yʇ5}4�V�{�b�4��mj��	��2�ҼHG���qYchSd��~��#��/�����,�z�)`��'
mQv���J�AZs�uO�ʢ;�3րY�έ�f>Jk�PȄw����a���x�<=���ע�{ú"���a��z�; ��mݝc�7��"��'ܟ�6�\��-�^�@8v�
�a!���^OP��3�		���{�����-�kJT� ���]�Q��!� g�9%�.�W��/L30"Z�q��tp5�(PT��R�{��������Ypy2V"?w4��Ī�a�W���.�CEb��#M*�����j+Y��i�����`baA�$��W%�Uy4/0�\��£�H��ܸOY�#x�����	��1��`~�a(�Z<6�u�E�.U[��&��	V	�b��NXY�$�͚��B;:��/�є71hx�&׾���>P��A�55_�t���Y�ǖQ��b��6��(��v-�w�ό��Y�C��v�;X�����e�~�'�r�.-���T���(��v��҅�e����U��2�	��s[-���$5s��h^�`��+�*A���yш�7���X��A�B�����
5��k>��r:<�����4����vd��s�\�q��EO����/��X��.q�ӫ�'p�i�}D�X �.���L���,v���&����7��(�[�9�]� �����W�f��~�@M���� ����1���fk6�n=��c$��1g����5S�ePV�����K�d���t�Zʫ�>����v�O?�T�
�"�"F���/���v32�o�K@z�8�yhd�mgK���Q�P\q�����G�� Ji���lD���`#G2����d�؇�z���Fc���
��h�z�"w��8��Mi�F�x��.��;����9�-R����.��G2���Ͻ�F|����M�l�}qĵ��c���{�𱻒S���ct�x����%*x�:��/��V�1�)썋���q�)��&�yH4���"<�u�hF�g�1���"A�m,����=� 
��5�j̦���^�B^Y ��\�pٽ��+���a��M�+�{�F����#��wN�B3�	��~޶qCZ�{�D��E���&���Uײ���3H��6.	8��rLE���ń�H���M�#"w��u�[ہ������@��l!�"�:�,��#�Qn�AG^��t�N�-�4�z/�L���4��{<�#9Ol�mK/�՘���̯5�<OO����J$�{۷z{b�����ɓAL���h�
\���w�\�+^����c� ~���@:�J&��h 	��
U��;��m� ɠ3���fP�/�ʍF�	�v�l�j��-�	v9�S���ɖ}�9��k__��C�uV[��N��c��rc�XD�~_�~��s��[?>W|⤓85.�%��gh�%H4{{�8��T�ԫ�48kU�P�F���*@�彃8?Q鿷�g��E�
C��T��ә���Q�(���8�AZ�L;T/��
�$r�7��\H�rOÑ�~��o"k�v	���1���瀅℥&xd�#T��š׭�_�D��%mT 2z٩�.x���9��rh����$Ӫ�Ӡ������r�Ӕ�Oލba�����}ę��v+>CMn�^}��j�?��g���U*�i*��U:|(%��Q_�:g�q|��}�w�v���G��1����W;l�^P/.���CR:��yN%�&��l�;��s��\Ai���%J�7j�%r��h'& j+���[D�j�)��CC�u��\c����
��,j�!�"�S�D���ʸ���'��+�����[i0kM؅�\�#���d�y�6�UP	�Y��r��mp�������^3�2Q,�N;I�1�|7�ј=���&Ӭ�i�!�n���;�HD[�j���xT`?���/`�h���*�����j�=��.Hm����E@"ѩ���ؒ��teQ��HmvT�|�8$m͇�T�tՐ�Y����B������������]�(��9lfc�q�$�*�=3�3��$P���8��#/�5�^t���UG�̗����Wғ_C��o��M���w�k��ry�a�3~�q&o3zg�9� ��[��x�z+q�:ݜ�S��%�r�ߪ?������'�C;A�C�=|k��������Y�YJ4Ei����Gr��vQ�CN��[�7Q)쥵��w0\���p��]��v��mr�O���Ɯ{J���ĴQ���z�mGv�Oǋ�6f1v�,�<�9�����C��F�%�U7\����{ȼ=bί����r{�ci�@X���-^&1��[E��w��[���57e"���jNC�N�7��m(��56�#����qG��%J6+.q�!�'y��*�	�Kw4蛒��� y$@���	9��|i���`���8�\�����(*�ᴀ�d^%IT�� �ŋ*�T:0�'c�":lI&�F$��Q�yZ8̤"�YMġ���Ų����*��|�3c�(}����C5�A�$�Ju�"�d�5Bˣ�/#rё����1�Hr���`L���e���MhW�5�2�k��e&_��뗓;�Y{j��� �B6��+n�톃��aA
p'1�/Z�W$�`ǭ�;�=��mi�_Z�љT�@i�t�aaHm�`�3��l����~����z��gB�H�Y	��.�nVGi�)�P��#^�j�a��1~��NY�X�|*�T7z-��*)�&>�a�� c�SB�_�Lb_�@��|�G�3Pva�p��y�6����(��х���p�#奬Sm��4�8�~��	~��Y�[����ו�8�` 'T͔�e��W>�`���I�$��T�n@��i"������	��RA�8֥�>f���^��rN�|9O�H�QL���\�h�{EYM���WO^@�O*�'�#	�B�h)L�	�fV��V�F%[u�m��"Ѱ1JmH�����s����@Zɖ;�ڽv�����]�w[����a����ۊ�� �n�I�!�)gWs��>�5nP���$(89N���+P��j����˅j�;�u�~�$N� ����{� ƺhSx
�CϜC�U�R�c�cB����J�ƢB4�z���o�D�H��m���փ��ol�E�sڀ�⭨�/��($X]�H۷|�9��V�`���Ox���6�������J�:�H��r�*gVtň˿�!W`}�A�bݥ a��HA._�Z��J|�[���=�'��(�G��Z��`j��<*N��&���m8��8������42���`'1��nM��3�6(P0X���-�W�0����z`,;�#V�}D!����f&W�9����5s�}���b���Y��-:�]!&{b2Gk}U�D]YpX�~]�q���n��Ρ
F���S�{hC��a4�m�����A����!��K�`���)Mj�@l[����]A� ;n�$��@��G�Q9�al��/�</y��z���}ԠΠ�������M���i�}G��"�E1���� 9M�Q<;���}���5b<�}��VE-Oc�� ~`�'(�@��=�����ߺ�?��]���TQ�ǔ�7���a0nA=S:��hd��"m
?��ߙ�\CXW�i����Z�4��]����C=~X ňW��������c��u��V�W�L&�'�F�e���(l��Yr���-%���?�.�����P>Z�N�Q�Uq��cD�d��Z�k�t�^;�=o����a ��`B����3��
���u_�����E3�qO�5Wy����ƾ�K\�K�:JQ���]��+S	�I�O�#�e�!5� %����ҋ�y�G;؂�w��Rd��m��{��Wz�&�#LZУ�ADU�T�Q����f?L;z�D�"_����ș�*�����EJ�a��M�|� ��!��n��"n�''�f*E�=��>�ar��A����P����FXTpԪ�L���"�4�#���P(ı�k����]�����{�t,zI�
�N��ȲA!���z،~	���|��h�x����)�5�uT�Fh xsq�����b�;��շ0H���<g� �|��	�0.�CU�1|�����@�10���b�͜���C�f�шG����v�J^��8^VScy�Ԥ�c���R��|�s����Q��)��yM+ğ0�p�A�!sF3z>��VUR���y�'\�\�;��g�L�^^m�a���������x:\9�s��]`;nn���E�Tx%�����v6��>���C�*r�1ڟ�V5y�H��0�K���a^�Odk���BxIrc�c
da�~����kM���5CJ|ɤ��#�v���QǴ�A�ܘ���QО��@)b���c8c�lՁ��z`�4q#���D�b�e����e^hN9ҩ���^�H�;F��WNݖ�6�>���J�	�ZT۩�:. <��7�֪&�+r!TM��#�'�&�ZF���ܜ�]3�ڀ��YN��꧁��yTiYBia}%DL���� ��9��n]tB0ߜ!6G�5��4������,G4l�f� �?���r�;{��#{jG~�g��d����6��?W�!߉&@���Q�d��MI�
��ܥZ�{����[�
h2d�L��	c ���C���ޜ�	�U_��_2����C`��7Ȳ|U��Wm� |�zu��'�]hQ�Bd������ƅ�䤝$��� YϞ��H���o��1��r|������r��r�4�{P��Ro�EƮ�xt'��C3��Z������EIdحȥ��sC����_�*n:D�Nu�7M3��4�8�����\/��#���;��q�Z~���PY�#hk�GO7��4 ��@ZNl�Q��	�=]iX9*����T��@-����^�ׂs����ԡF��v6�(�޴�!���wm�h�A�)eE�:o:c���uD]�/� �N�9���wW�X\:z�8��0*�T��.��.��LT`�pz5Vl��X�P�HݡV?"a����Tk)>����f^�p����ar�t�������D�uB��u�<\�V�
ef���/�l>Tu2˵'�2<]�2z9|�p�� �b��a���4(���՗Wh|�K�J:(��`��^g�_��j�AW?,�~�J�Q�-gn�p��Q�?�7��wP��( ��1j7Jӣ.5n�����h�A��54 .�&*"��[H��*�� �ޛ*T���N�	���tR�n�>�諱��6a�V|�q���J����Ӻ}xB��aݯ�_o*s?� �og�ߍy�%��e5@�1µ� [e`��C g�#c�uh�|!a������
n��mW�<�P�٣/��>d�9B��Q�^8	�V���?��ǂ�����D�q [����R`��Z,W��w+��a�e�2������'���\�C���j|����OW ��3�q�ÙEn�SY9NAr�j=�:L<�-��.I�;�H_��J��U+���G��XtM��5	�,��<i����S�q3���&��8Sit�H*X��9j���$����Q��|Ib�[@jL�vC74�X 崂����2퓡�a�X}|�i��͖@[>ѥ�g:c�;���V��[
d9I*���O��mԶ�[T����+9�KHf�~@7�i{���*l���U�6�q�~��B,� M"1� iA��]���X^
H
�^�I��ฺD�Q��v��t��=rC�5h��#� �4	畞V^ ����I�������͇iJ��<�˴�,Y�J�KB���`�4G�ډ"��*,4����Ij������4+&��b,v^�X�9_�@����тg���5��i;�^8snH�K��d�a���m�Qa{��Y�1A�� /�ep�zx~c?"�����:`ua��\��68�a��֏�G�Ff����'����C�0 ���o�ogO�e75��O�txaw_�7����Wߥ�V����1��?#p��9�q�9���C�k���E�eQS��X�^����G���0��nK�=������F��]�(�ŅaZ>Λ9K�K�ir�[���d�[�K���M]�9N�m�����x�naN�u���0u'��(��;G��W��"�����V�����qH�m�1�t���M(nƉC��ck�Dw�|8}�����DO�P1(3��˹@c##�+:����� c��F}��=�\���.K/�w��]�����a��I>���.w{�-�`�/���%���,\�^d;|�K;��}�tx�x �������(��޹�A�f�*�`�W�G@�xE�0XJ�j���� ������\�!��}��`�yr\xI"�	��E�DIȞ y���ԟ�{����,�Ԛ�Q1��(V�����\*\hd���C)��AY��l����8����ѩ&;�U֢(��K�R��/��~I�'���qʄ�bջ�����-J�!�dX ��h�$�%̸�_�űr�[!��
[�]Ah�FG�[R��|��^���*o�2��p�6�_�o�?����-̒ �6vf+ش䎢���~S8�v浾@ᕂ��2��Xaiߖ�ѳ�>I&51�����nj������� �ml�6�5 dR�E. e������5V�r�"���!&�@`��2��g��Q.m��X@���n�6��"ȅ��>Ś2@[#�;��Y�ѭ�����l��y�O��XN���U�~��>֭1)�^M`���^0��>���6�x*���ڈ������"�#�yB9�]����K0�%y�1ze+�!]>���oͼ'tP�z���Wtq��=�,���B�ut��Õ��e4��g��Ղ�~_�9b�/x�KO�XnEk#�bJvO|~L ;�����;H4�6�S�ӹ���|GQ�,���A`�ҍ��9��\�����M~ v����oPr�Z����z�5j2R��
�U���/U�s�'�&:����j;�[��d�$S>�wn�kq������l�?�/����� |�>Y|d��?u>����^Rv�2�v֗��26��凇S,���"�5��/��I]uX����sV�OG/-݉� ѧ� `�-a��.���h��C����dm��;,��,0-=c�_9����S8�ҋ�w
C2?�f^�`�da<�����4/�4�'o�]����,��gj4�� f�B���i��D������7�j�+&e�z(��X"������s�!�W7�E��B�a"�j�x�(|lH�&�X�.�׺}x.��EZ}�Ul���6E�rV����_�4%�y��6b�>�5�N>ҿ��	�0B�ly�c[p/=���S�~Oϒ53�@r1�%�ޟ�ˋo����
}��:/����E\�Q^~�Y����a5)սtȒL���̡>��������Q^R[t��x�8Ӹ��\�v�`׭0��"t��6s�^���E��J���+(A���};X�:Ӿ�`�U 3%��o�ʚ���*��̡b�i&����,L���<h �th��ҏ����![���ז�V(��y1^�rOIx3�	�Eɕ
�;�.g�]���L�.���c�?�υ%�1E��
�a�h
��P�u]M�Z�`�J������֎��f�_vW�X!�1o/�C&�݃����|�,i�E�L�� �Z3Z��Pi��ccV	�|����+ �q��=͝W���|R�/2��+���`{���k0(D��WF�~%����8�����<��ͮ�GF�7�-�|���I�!��=6�&��ܦv4�d�/<*�Gͺk;��p��TT��&�ם���-��l!�M�d������o1���3H�_Z�B<�n׉�ZZ�����:o��MʗV�*H�X�9(��{z|7���͗e�}6���tH�j(�-#����z��,nX�Ye��K*쌆q:TW�a��k�yA��25��#NG�����D���F�F9BM������D|]8�ȷ�5K@k���s+&�A7W@R]�o��n��_�
�l I%*�&K�
l	w��F��̶�\c-���2���?��o�֕՘`ثF���uZ^;+(��6ɶcyG�9YQL�#�o#��an�Xwn�ht�
�H��_P���r.q������?b��Y�a&Ɉ�>
['X�G]���-oR�y6���0�&sd� UP�t�'e������)�|h���c��v����ªj��g��\�5�������S��!��=�_�jޔ��}��Pc�eOS�P�A4b�������|�v�z��^�}�lZ�^��ߖ"��!o]k.	kvU2��Q�cg_(�.A�KϏ����n�7�e��.���>�
�Y�Kq�N��ǁLhł�i���|̡��h{�9��e���ܥ��ꩦZ�6�"�m\��h�|*Q�l�*�����=����c�+e��,�:+LS}�\C�(D.K��=5%�,�tܛ۟N|�DѤ�s�>i0�K_�%�3�}^���"�7nײ�J�����@���%����m*i�&{�٠XǍV9�ԇ�%И��$��7\��fb	�K��* �j����+����/EW���ѐ��5��X>�m(c�%oZ�a��� ��,t
���j��x���_�N�DV/���m؁�����6��h�������G�.KpQ`�<�R���v�z��d2=��?Y�T���z/���@����hi��\^*hO�yW��X��)��8�`J'��vu5u!�+"o>S����@Z�T�9���J�L�}-A;f
���ܭ��Yױ)f��61�dyW�K����i��~&Yl�F�Q��f .���ׅ<Vjڻ4��V&��"B��^  �epT���/0Q[�r?B	kSV ��}�W���K�J&��#����Y4gF]�P#���o���9Ӏ`
�K�X�w����y�껇>�c�=��\?m]\�b������8�����,����=Hż!������jvkA!�/ii	��"Y,4����9i�mq�ᤐЏ�D;w��ͅmTXs~��u�vm9�� ��'�������E1�\i��]a�dLo��De�	��`��0%�7��]y���C�:*2-��=f�'yw�"�2���0O��f�ݧCx�e)����>�%��򂵰R]�
o��Zuy9��G��૖M[�Fl��� �rGv=��hW�����<�!i�`
x�݉�r��knX
��FE$BS�ν�i删T+�Cv3J��F��
jl_m����	�(b@����v��TAF���	?�٦�"��u�����y*68�hE�/�<����Spe�9�6�b�['j_���F<0�J�'�r��*��4�Q�Q;{k,C����S��`�^a�|�a��
o �|�f���d>�d\�K�Ծ��!Vfy���k@~޽�Kٰ�Ala�T� �@���`RS��!�<>蓫O�6�}�o	"�=� �?��[�����I�o��@����������㸣VT�B�������4`���ȫ.��Ӄ���EgM�yi4�̂�4����a�:t�4��K}��'O�5�FŜ+t�E#5��=�]U��0Ϭ>�;����$�۔��霏���D�N&%�m��2�)v`���|Y-�BO�rh���Ѵ�������}R�O�wl�;%:�j���/A��N.��'=���<"b�j怘�7?���o�i(��4��	|�
�eW�s*7�^���}_]�[��_�9'�r�vS��6j֞�9�Nu]�"*�+�>��5(�����Z��@�e�)���@s��`�
����إ�{c5+��(&S�w�R�K����>f�k�`��M��2X yd���Wo�'�7��P٨㫲���q�<�5��B�"H� ���x'-��c"��5A}�*�"ӻ��3R_6b����2L-�4�9O�x�|K���.roa�~TF,���yyd���0�z�'���hi����?qE��P3^�wJQ�a�d|��f;p��,��ȷ���#[�𰣁�r�.�O��㎝�-�~�X��qt=�����Gd����K���F��H0�rRX�-�3�M�?�RR�j���s����쇎H��Q�`�^�p_^02�I�[��A���.��8�H�Q���a�%�U�ٴh�x}M�y�J�[]��J��X톨Ƚ�p�]&kJ���Qj4�f��)BD�e���Ծ$Q�CZRJ��[$"�7�M��й�l�\=��,A:黨q��R?o}-<dFI�!��g��˂}lU�h3o.c�D�7[��}����+���r=���hIV��#lh�fLQQ��Pt��a�!�NA/I��I���&���D(��\@��e� c5*<E��4Yq�i�[�̢>9M���~7(�;�'XD����̘��&|�R��˛(�f3�{�UC��&������o��i�ө�6=���v��P<�W-����?�~��ׅ��Q�� ���!S��5��4Ml�}2>F�2��s�k�]j��l�Ɠ�~K����5g�iTF�Y
����H��IUd	��c��c�����tјX_��so%P�o�1'1��ᯬ�����Xr�a�?V
�i�T�ɪ���W���7F��4�sos)�e�27)hk��[JRJ���,�eBX�i~iF`���W�����\�^2D��LW��p��\:
��O���g�	nf"dÑ�
'?f�I+�	�A�����>���A<S������lh�,k���2����-޹��hz�!��/��=LYa+�l�F�6�,��B�a��`*�v@+�`����t&'�u2�>{ LEN$!o1�7Bzߵd]�c�}:|��v�-��(�t���k%��iQ�R�$=�f�~�%�'�}^l���4��[��ȟw�T����55�<�#Y��/��ݴ>[�'N��A��׉#�}����5��@��}�o��+�#'�u�>��+j��y� HD��HL��5�a���Ux)
�d/���3��\=l[�	J%\8���y�)���>�I�_<��O�R.5���p4�0��R����QxGĞ��9�r��G�@�9s\��7'��c�2	>x)E �h��Z&�����q:[������lx��� 3�S�ͱ��0YCob�	=�1zqT�F��h���b[%Iٻ�b�-�X��מ�al���G������8Ǒ��UQƁ���D-0[g�Bu�bFZBۀU-�X�]'ݕ��%!�c���U_�j+8�Ӂ-pĭo�W~!_���Ӂ��-#_��ō�˓���1k�[�m'�Z�ɋ_W��{�mzY��- �~�_���x��z%}{������<����ք�L���S�� Tpi�x�xj��	`�I�͠;�>�: [�X��0ق�J�S�N�̐*�V��
�'�\�B� ��>�a�?�Q�ա�x 9=�x�2��έe�DƜ��o��,�=@������Vw�k��2{���n�_v��<�Y �o�����!�!H���;�P�� �19�w8�9[F�R���^OA�F߿kL���,�������g�����p���̊6�T���8M�#���Gwf�hg��4����ꘖ|J�6d�U &5�~&���tYþ�RP2��y��Dȇ"9/�D˕;� ���L�Q�n[��f�D���Bo��=����T<�&2�Ey��%���D�>�(�!}g���/X�`$�-�M@uf���DL2b/����`���a�f����K�\�z9K���9��S�|�(���=Ջ R�y��+�Р_�T�e��y!M�XLI>M���Ȧ_�3Y���+�7�U{ϊ� �r�JqF��e����p?<J=�K5�I�X$�������M`��	�lp|��|��ʅ�_֧8�L��fϳԀ$�ϣ��uѝ�LV�|��O�t�q�v�>m9+�3�w�kѬ�6=M*�j���}��vD��E�E�ĉ�MuA�=��J,��e9��
GT�B3�؄1���?"J<T; .�:���l�"���c��x�&a�e����42�A�|�'�u���ԑ,��D� �+b�7�-���^lw}E���_;sa���@0�x��%ol����F*�*��^|��np��ZK�(7g�u�^�����*P��P(ۃMu��1f6��~]��#��������@��EL��[���k��>q'x@�i/��Թ�O�O�<]�3#ofp�,r$녜6��T��:�8��rX@�OZ���A�)�� �s��2���2C�,7�S��-`������f��Ґ��w�f���m5No�x�0�E��VzU�k�G�<�4[��!x}���磭�CRǽ��q�1�����~��8�����F�)�8t�4i0#��g^=�H��'����7�$(��"��,����8�2f�(�r���a�"_^�ۘ*�~���=����r�F�w�vk��?!������fa(���+���ܯ�?�E�� �E�	��	��#!��-[�?H���l0'Q��%0�c�D�^96�Q\�a~:�����,d۩��(i�װ�ļcP\�������ü�2C��d���}�W�"��4��N�}�_k�m�npR�k�J3�eII�g�J��kK\��E����v�����Gi�4b+c��^2ڬfO��7�!A�}\�ֻ�X�(����*^�Y��|��������n����*���\3ɾxF���i[��$���C� f��b���������J��s�%��RVZer�h�niz|����j$�u�*pi�P����g� I���i:�nK�db���"���`U����K��[�K	li��\1�7�}YA.�#����B�6Κ�3� G�O*���ϛ��'�"��_�xB��!2w�`a�yR<�~�+8�1Kzԡ�\.�\
�ݕިj�����M���d�һ�E�O�=3��A���~���}��u��h�� AФ��L���+ﶶ��8����}���gn�Z�PC�IU��[6���12�}^a�2����nfi�dgtmQt87��`^{�pz�Հ��1���r!]`)�ØHvMB��iK]R�մ�!`�������eE�Cw��;�:�X��Y>��~�z/�6�Rc�>,K���1ad�*�S1������-D��������z��)��N���1�~�j��͉f��@kF����ͩ�5���'4Q��쏌��]�$� GC͖��y� ���k����;̟�K3P��
(j3:����*Uv��1�?spD��Ž�>8��]/m��Rb�����m0i�޽c�pR ���]2V�O��|2��yṓ��-g�HǠ+,�'��C�Y�����a��b0��ޔ�͂���d�� �!�,=R)o�$R�ͼ�N`�������:ٖ,_�U��
��1��ߕ����+�i�V�=��5����'5�)��ѭ�����͢�*���ҧ�Ii��(��=�,3�
(:�W#YO�-��vŵ��.��1�g�_��ZDDǇ��&��3:��L,.r���d��h,�Fs��Z���Bo'§bd՝�]<�,!�~�^���5ǚ�{�#�0e��.����KB�I}��nu�֬�M�ƾ���%���x:�}�9
�6��&���0��#��+t�s[Y��8�4��2&RUT@�R�\�6�貣Fo�$�P�D��{��ͩ�=�tW�i�g���ɦ���RA���(�=����Xw�%[��um�M�z+c�N!��Su������Y�3�`��/g����ӝ�uA�b(�l���N�"���n����]��CX΁�n�@Nu�K:�;r��b��*D��ic1kM�q�E�\�1l1�� �l8��<몧�'p	�����Ni�t*��e�"+ ���l�/rvb�����sX��j�jSi#0��>��H�H0U5#�e҈�b �#�
��l�'fm���ʹ[X�GE��Bؿ���k��y)I߷�%S �'{�n*�)���*�k�FH�I�cYdR�1fA���tf��1(�&5�fO�؎��AL���3�ƌ{�X��ȱ!��i�(��$4��֪_�\��r#Q_@�m��m��b�C@��$Cp�~(�~Hup�R�[��`5�M�&{���ZlWC��d��\�¯���Q,��J����*�E$Q�<���CtRv�����yt.F0�.+ 4�؂��g�����i�	N�*��wc�a��:��`	��G,H�8���>�<�//A<'T������uh��k�M���/F�o1�!�="6O%0�I��Ʋ�ު��g�u� �g������/��$��u(U&&`{权���7,y��Y��a�.�Vq��QB�Z�5�;iZ���@��V��9&�1�� ��w����)0"��R�@JzW���3�<4A?�l%��.l��!�X�e��3��%���
S"��]М��H1e��c�NF%�;�	��=�M��7[�ܣ+�����(Ɗi}�%�C`Q�Pe��<�mjT��Ԡ�G�M����b���,�U�!7-�ht}�%���:ڌFȷE�Y=��Y�@a�	��`��D��y��������&g�}��M��+M�ʤZ��!�4���a(����V�LxM<_݈^�;=�Hj�`)�rr�� ���.XQ��Zp��`�v��NC�Eƻq8��4��� ��@��L�x����꼱�K���5�e��]���}�@rG�6��Z����tv�	��0,ɕDD/�*tQ����.�����f�^FL��(�tpD�&)R���\[49]��V�ۑ8��u��̬/�
y���o�8)6\�Y���*��t�^["�-�.���U�PT<���2X�厠Q��G\Gt������ͷ60�n�	�fiU��.��n����{g5�+����D���Hzgʠ�5�I��m*��\G���c�%�|]�(n
�=�U�D�|A(���9�`a_J�WaMzNxA��3�Ř(�����9^��c~�K#
�s<o��9�X�t��%{l��⣠���J5Pm�cs{���\�'�6�#��CoD����*���������8o���ȑ��&��D\�t��͠>�5�ܡL=�i�8Vڔ���J^��l���$��ƽ���)�f���E��t���q�>F�O)�p��X�R<W`2��#]��Y�:�=R�Xq�d>�3`w��A��� I/�$Az��;�@���|����x�||6`Ӧ|�;��`��!D�l�>���X@✱�I�	��俷+}3ٍ�ʅ���'����ٲ%�,+���u�$� ��ɩ��/����G�d�}�z�8��o��{����GeH2e�?ͰS��f���C#q,	��)�����l@Wt��|hw�ԋ�*�~b }O��E���Ի���'-/+���/�+-�~d�s�ṣ��h�L'�<�Zτ�]�����!�?�lDA�CU{�HRi���$�ܦ��p;D�2�EUC�*9�������E֐�Q���ƴ�&������zF����I/=	��&��(��������x��P=雏�>���N^�r��4�ys��3N���`���Q*�22�r�Ӳy ;�h`9��U���Ib�{�D�di�ʂ���)�r�E8�bON���v��:,�*�鈝?�5ͦ�j/��/��!Ղ�Y�\�c� ����GF���sn,���~�X���w�I]�H!��ۨ��2k��f\Ǟ@�8T��7H�����e�9�"��1�����t�2����/5�3�d?!�՗��R��C�l��+ف�����W�J�x\#�����+�k�bhf����)�H(B��L�8QUPA�B8>8�dt�k"��cd4߲^����)n�1w�M ��,���f+!�a_߿à�,� 1���لe�듷��1=���.� s�eG��t-�b��vs-�t���w�����c��UO�;���w��55�3��pa�ޞC��-)�ð�r�?��@�,Ń)ץn�}B�����rI,���5�t����H;cS���6�d�k���p�t���|��J��v,۽ d��������#�v奎�:�J��ɮ�j%�_��M �Œ6�ZQ���M�2���W��Pq͋��نa��,�$t��!�c�:��y��U��za�>�N�����U��N�>��$��/U��^p����S>K��Tǜ�����j��l�������Ӟa�09���1S߄,>#���x�3� �q��s��=;��j�ÿ�2%y��:eq$j��SǪ�}�16OpHt�>R �~!�==
��8�����oA#��0Q�п��/J����V��^�c5�A�:�q�tEW��yJZ�ʑk�^�I# �9DS/VȲ�������6��XO&���P���5hڽKm�vkMx;�!Q{�L�hk]�ãa���f��M�X��I������VofzWq����
��<�^���O�x���Y����J�&�ٓp���lV72b�����lMi��7���
�%b�.񲒅����(��q�+V���>���.Z`M`��������U�y/�Ԟ�ٟ����tY���s);��Ļݷ��O��̈́����D�������:�%�:�v�|�@f|km�q|����dF����oɕ���W{��tz�{�C V
�H�\�SN�u����H۰����<��Q8����:��u�:�������o����v��,�B�w��|�n�]�(j�+�|���:j1ǆ���ubML��
�j<1l�S��	�!�d�W�\�V��}j�I�y�R�?/<4a��_�kM����A~�n]�87��'��z��n��PP^��e�	c��R�(�9s�A�� z|�02IÑ��A	� ���?5����U��r��1 �ND�։7:Y�L��s�%]Pͩ�e{��E&������If�V��X>��!M(w n�c֮˜������u�h�eK���>q�G�R�E���1*��"���-@-�ӯ�����+u�۰����DI�&�u/	,�3�ooВ,�*LA�ܳ`Ώ�|H���|c�X��X��K�+ ���a!�$��KQ\]\;ؕ�o2@c�p�k�ig�!�x���a��5:���y!֎�oKt�+ ���L��I�ҷ����?�?�d*���Ee5d/���P�L���������Nc��/`��$�$���Y;-s9#AC�y ��<w��'�hA��bo�Dpo�v��;������zZ�<�nY_�Ԯ.Ѧc_[V�X�hWH���U�&�" ��E�l��S������ �=��Y:4�bs���%��9W'�|���^�ސ!|wU����VJ�?s��3�̸�h���T��1��Y�#�8M`My����D��!"�W��iG.-�e1������mzswZ���6�x�t޿P�o��8Y���ᣗ�]ТN����FH�SVʦX�4� _�����';ts�b���Dw�����ݒ��S�6�P�� xF�s�&y����J�5g�0'c�u�9<̠Q�?;��0�tP���\���0b�<����	|�H~��������X*���;��?V?�$�Fſ�˽�J8� ��̊J:n�./�w���N���Q5�&���ǌ��CrK�����wYJ�r+$\���vy� � ��,��-{`�}�+�]u���77#^�a�)Dt��A�d��^U&\!$OR��P����/��%�'cI�+֋��c��L�J.ֺ~��Ӟ�X�y$�Ib1�!�:H~�
��8��_�	���$��F�{b��d��u�|��y�M�,�QZ9;���W5I� J?�p���no�#��]���G���-پ�gD�\�TJ�'�4�>R�	b�G�b������LG(ȝ��I����Fp��OJ{M���+
KfgvLW�
��p=�֬:n��<M�hn	�&ܪ�Gy��N�t6s�c.p8`d�~������HMvY������!q�e��.�!���u�19H��k�C��������)���F���	�3�l���x�l�cj�����)�R@愚Y`�l_`�Ԡq���-պ>�j�m2�L�\�[����b +����2��i��f=�x�0ߊ��<�Y+���?�� ���/�u�K����+�G
e���	���9D�Fʺ�t����F�vKE0pC�Ah�Q��'J�Qu:M>wך���G�*�E t13�?^�z�i.	{���5����H��1��1vs���z��(�΁�B'&�%VXl���xI�DiK2�_N������S�����@X!�_��(�X�7�&��`)\u!vȘU�6<�mU�ߺ&����
�7j�m�	� ���Я�)y������D��Q��p���P>W5PS 4�U���_���c�|C�ECN��+��u�C8籭f�m�	�Pd4 8���� 9T�Qp�l�x9m�m�Aȁ0����.a�q�<ji�P58��Z���Ԧ��΁v[ۛn�4+.�]�Q����m�]<�N��YN���[LB�8tJmt[�E���_��Ex�3t_d3!��'$�&�g�F�Pe2��hWl��ȯ�b����yҽ~j ��MLE�75[�{B���$X,�z�nkh-��#��	� =�;���hO�IJ]���Y�?��Qn�Pe����.�����S��9�@n�NK����T�-4&p�I˶w��<�\�:�h��^R]�1 �����ݵ�4���?m{�3-�Y"�:!8�;�e�6��}Y-�郢�C�{)�z`���Ϫ���/D���_���1X/2���L���Ub[(q
#�UzZ� ���P.!��K�R��=�Ĥ����[`��\w�W�9P!�ӳ�e���V�d��*�k�Y[X.a�ȘWG���A��Ƞ
b<E�5a7F@�T⌏�e�W1[�$�D%�
�u�I�J*�Yh��th�@q��b�����8
���t&Tt%X3Ъ9m�ͽLa�ג�[���K!���	+]�zI�����"�Qܜ���y%���sI��=�h���jlD�N�k���[�5ڊd��;
�@c��:=r�~��޾���po	�D /ak;�Iɉl3�w��]�s�&�z2l1!N�c�Ѳ��R�z�Q�7Zi��
���M�Pen� >�����D&
dq4���+a�f�������<GA����
j�@6�=�Y��k |��Պh�{�@����.o! �FR��ߥ<���ٙ1-ҋ8�?�|L>-����	6 �3�np��S�����g���bb�Dr^*`o>e@)��ja�<
l����m�+��/[@|(��{bP԰&��C^tI��My�b�����(�^��B��:6d8ŷQ�ݛ�96���HB&�.�����`�÷�3�!VQ�[��)d9��]{�����u�6~���Rm�)��--�_T�sV��m]�=w�U{��n9�/�jޔQ�Tf�2i�m�Ō��y�VQ��5����A�-W�se���+6�(a�߂����A� Fˆ�R�� �h�b܈�`����Xl��,�*�0�sh-�
�'~���5�&:��q����P9<|��k���;hW���22���e#\�͇¹��+�@�ZRcN]�:]��Mk0�2����\Z?��U%���4䀑H�2�n��'a8>9�Q��.rjBN��v�����/�SHY'י�4p�yĖ�,��lM �C��Ő]���2F��G�䁛�9��*Vd�� S������Q��m�n2���ɽz�w���/h�	�,DԼ
o�d������BG�dbf���wI��F����a	��(�Uu> +�~��J��n��m�'F��8,k�iRy���{̣?�X^j"H��&(ހ�ó�ǭL;�iv-˰
x-�P�9"�c.�pzc2����`X~[��p!�1��3V���$�30Q�������!�i	,������2�طaHy�e��o����w�:����A������A�{�E�MNtǱ�xf�����u�j�	
I`��@@��æp���h�"�S���t��( �7��m<#�ǰ�`7z���N��<:�Y=|�֮wɞ݈�om���7r�ܧ�܂Y� ��ݳ,M����9�ُ±ϰA�\�,;�K�NT"��]�E�ʣ�dr���<��*��P����㯉w�A,�pQ"mL&�,��	iUa���TQ�؛L`4\ѻ��E�v3�f+�#�ԓq헪�uv�
�Ƨ�VCK�Z<E��Z!�i7IrHC�9+���(��%P���
�hLł�A�q{K���(�fO&��0�[��UԢ�,��2��̗tˆ���GYt��Bso@A��mOˠ���d8C�?���1s�j(lg�6���G\�����ErA����Q��̣@܉5e��8w�c�����N��hZ�4�F�x=Լ#�ϼ�R��4��ѕ}Ŋ����$#5D�a����H�=,�k9	<�+���|@���M��n�w�/��Ɠu._��9��a���N�`�`��cp�I�!8k�*���Ӥ\��o讦��:�^�O����/��XQ&07��)#��Z�_g�Ep�5��C���G����C���/� ��rZ�Z��l� ��,���^��KTJ6K��ː��7��Z�IF����6�����(�x���~�2�$P�ud��#̊8�Q.�D���Ԇ�Y��M%*m��Bk��D�0�9W?�C�*D��w���D��j-6����8���*����DAB�k^clM�J��Ur����G�BQ�ǹ��3�e(+�(��%y�� Ӽ��ާs�]���zC�]��Ľn�?dP6Qx�v�||��CFt҄z#v\�etʄJj|��`�FJ�{��KK��)$շ�^���wDx��tl��  hҢ����8S�������qY�g�h`j�ڦ��X��l�����
���'� �O��}���o�hY�t��0WE�M�ZE nZ�G���Ӻ����JO�X��Y�a"8�+��"-�װ
��?#�������Ř[�ђ�j�r�����R�zEf<���1S�YʭNs����4���_��=��νˊG_x�ۼ�훼����7h2هĂ��Q*�rOd��[���D0��i6"h&�$�3���7����  �7�a8��Kc�D"=�j9��C�C��1�,�zV�jma0a$�����$&�����Lɐ��L�?ӑ���Dj,�:6���Bsql�n�qV3O�,��� �@����C2�5�F���ޖz�YyskE�_P�a)�a���<�S�WP�V����ncC�b"΁�i��>����usT���a7��Y�;�F�A�ަ�FzC���5ܻ��</�Uw���v���]��@7H�@3e�s$�4
)���CDq���� 2�&�E�9��?'��dTd}@��A����uu.��G�/���Bj۷�v�?�r5/��ٻ�`>绚C�\,�[�c�y�t��a�%�ʆ�$�z��*F(W#SK�$5�1�n����z��|��`��w2BL�Ȇ^�1?G�A��iN�f)V���ʻ���h�����6P�xo�K	���F�M�=��/�@3	󧀀�q��m9���R���F���m���!�?�i�X��d����~��$�8Y�Ja��|��3E{��MH;� a�Wڻ�a�\{��x8E	`�kpF�
(����a�� ����0������ԛ�1'�b��c���f�ofh��Ae�޻[!�[�&���i�u�5zX�D����c6��N�~,�(zL8��*�b���R��m^3K��{�N�۟� �]�b�O6�j�eֵ?]ǩ��ww#Xڇ��D�[J���o�G��⋕�F!E�fA�I�n��^�8�s��V�p7��A�n4n�#IV! �q1mo�������t�L�~xk�o�J�����k+(M�3�5:�˃��X���X���zz,�}�S�҂��ʑ��ԻU謟�#U8U���.���h�,�2�
���T�fߏ�S�"?���òr�VCaX��W�Rx�&�����I!�*�>>����dHK��9r����;�x!��/p&�G�F������c��`3��&��cq��;U:�.b.��Y�;���ZF�H,僙'���Ӌz�+�g�*R���g.4XWA7���+M,���"?)c�nM��uvS� �A��,ͥ�)$�/��{,m���ߴnL������u��|:�U�`������H�n��)l��P�j��TDrR�Y)2��mv+��
�#$�ꉈ/��M0�^3��S�CO:�Y��Ԗ2_�F��H�t:/{�r�2�Ej���:�w5���������L�~0F_6s��AiT�=���U�l��2!��-|��gHI��aa�8&=�qD���.�^��y>�PT�,��9���^�85��ۀ����8w�����_���N�_t�:�����#�����@�n� S���l�4����sK����<Ƣ$=���	��mU���ӑ��3Ҥ"�?b�8����̑.��x����x��U�O��׷�=^H���kԊV��̟6����!�~	 ���b9�y[5�$vΞsX|^.�0��L����B�����髈(Lu�PnR�!߈�<�K��j�k��3��tâ-A��q��f��
H��?��ՇɤUE��,&��qq͹�x����G1a/�r�!��P���a�+��O���;�(�)|l��1�R�NK �ë�x��_���[o��֤�Cg��C�/x���X�b����'�J-�<��k�^��4��%���Ǎ��>8�� �E$B�'�3?v���F����Fkة쾨*�k!�� �+��t�D-��R�r]������<�Z��la|�ϼ_�Ɯf(���,�6�Y"���zx�
&|�\��h�`�Ny.��7ڲ����^u%���S-X�?�S�C��ngg�O@9�c��� O�!�BE��n�W���M�
��G���u����~�T��z����ׂE����p?��I��cP�+�;�ŗv`Uvk�f�u���GK��V��A5}����Zz��p^s��;� 6s��F����?�bo�C�T�FzR�qx�����P�r�ZS̞*s-h7c�6��@��p!0"��6�˕�Ռ���(j�/k8��?�2���
xa�epç����r���Z>6�"w(`����S��K�w��$:�5��c����3�+cA��M@מ��O�ӧ5��+`�|Jٽ
������X�y�0w�r�:'���*�0�e~ikނ�a!?Zs
��١�=ՙ)�:^�li�ƹ1�t���WTVF�� U{fnA��lo9��5�y�ƍԹo���.�����o�m^��)
�-�p��L��+�c<���k��F�A/T���)PxE���Ǣ�3��³�WM�����:,	�*�M�Y2J��d�F�bw��fȸ+�e=�]�u�?s�w�[�C¸��� &/�q�~�����0�b�]�a���+*��*�1t�(4J�����S�����5՗Z�fj�_>��i%��b��g��,��CWRIsB�\+����5�L2X4�')Wן����y5�Eу���+��lS�����}�\�	+�6�0��Ȏ*r�Xǐ[iѠb��kʠU~*Լ��[�=��}�`���Vq�ce6�Ѫэ����/�.O@`�T<����i�Nm���E��tBP&���1�� �?�Q�A�J)��h�I���^h�6�����E%U&��OYX�6v�a��t9z�LTr�Y�sY!���w+5�r(E�\a�9̄Y� �D��9������9h�HG�H!f}ݔEx&x��'k��4;��γ���Uf?ȝ�ON���ǨX]A*5��P8�B����e�Z5�=�`���W<K8>�x�yR[<���ˆ	!߀Ze�L�=����b������Z����XSUU!F�"�~u��z2&y4oYQVD��YM=�.ߡ����	ǜjm�z.���2����T�o��2�=D��p�R�:��آ��g�)t,���<��h��
�b�F{νCbJM��]�)V��,�6x�Yn�`룿N1	�Ҙ��8���F�^^�\_l�$�L%�ߥ9��
�az�²SL18Q!��?�w 8��z���qE�<���P�D*��`��+�E�7��@�.M]Y	U���9���GZ.o��L�z�b�H:����*`N�� OBXdv��1������ۃжJ�ҡW���2�r�2(,bn�y(��������aK�-�c����y_�E76�m�	��"\�_�
dK[���/�m,|r&���|n'+��������肾oD�CK�G�<�Lz�1���%��<��2M�������<�сۢl��Z������-����ixSl��{��+����r9�
P�]ԣP�r�ZR�7Ƥ�O)��@�[9&\�櫮5�ЕX�r��<�w�׉+q���j�51>�O�����0�����~. 1E��_1��Ы�1��`^���
s+8��Z�޵鹫>7	��:�p��0"�Z2��8'×�!��D���	z��hK��=�,��N=U��q}F�?���F!��t/���!��̊ �j�k}Ih�,Lkv����8�g��>����vG�t`a+�f%v�mgz_����F�(Z��=Ҡ��v�LE�VAR��Z��S�!r-�M9g un��?%��;|�<��f�x�(=|&� _<�mI��FI��������ʾ]D��Y�J�=�[��rn���?[Ɔ����)=��C��Jj�fĆ�Q���^[�,�f��=4������h�5�WG��=>�a�\0('�k �pޝ0�!��3����,Q�׉QoN�T�h�g+��j�By*��H�-W�6aI1��4�	�ItD�֡A�{�$Q���e��&���#o3'c���>��t(���|�OL N���y�+�8�fQ	0��|�-no�!QK���o��Ak��oK�^���tJ�4}�"��Lϕ�(�	d���2r��g��;��2��NKI"��Q�@����P�o�.����a�XEe�A�4�EۼG3!X���� �r̍yKdw<D�Rk7N�R!����ۉ�YhD����|;6K��2��X++���.����l�/�.�O_�C�j�q�Z%���[Z�?�MoaI׻�wz����ݴ��S���XeFǼ 'k�|qTHg%�c�	�*M�����Yr�e��v`bvv�,�h�I�p�80p�PL�h!��:���*���I����1�s��(�w?�jgke�T-��������Fߎ}�.|~h�h�}�*��i�)��I��Dh�!�!»�(�2/3���B��\D	��-3�0�zd�ݗ����m���s�)�Y5u#��?M����bGo3�D��t��u��_#S^��E��ܤ]�QE��J�%���T#.��}�~��p���8�}�I\�FoJ�%��Dʜ
����؜���ݻ#�1�\=��4;�( F ,�͆�4���%Ԛ��_�B5�B5�1��s�8����#ʟi��c�ڧ��19�/8O)l]n�Hv<bQ���>ⵖuH�|��~~^�B��Z�>[]��e��X_� (@�
^&���Oo
��D����ҽ��_�2mM����&�;�7�����&{�3�x�P���`y��iӤ1īތ�h QMd�n�-��X+��o;?-�2���5��Y�hK]���p����e��l,}L�}�S�:�k<m�R���؁�E< �P���imgz����h3���+�Ջ>�1��Y��my��pWf7ͤ&���d�f!/Ӆ⭾8aY�(����%~�y/	)MNy�7e�o�c�d_��9$�OD������HGve	�a ��1�(�Ӈ; �$����Ÿ㟊=.�PY�R��e����B���(�"���X����s(v1[o��~��L�B+^�v���x�D$�@<b(�y�m�4ξ0�\��x�r��e�oМ�9�����r��|oV{<�U�L7��FVE�fH�T��;��x�u^�d��t>%k{�NT�Ah��8NcZW��9Q�U-�~
���%@đ�i���q��M1븬�p���I�N���<���:��ڱ1��&O�V���(�@h�Z��7�m1o�ћ �����H��G&񢁵#E{�Ƣ�Dg�/��'�U'%��]�,&�����5�.��-��s�؎.�ц͊2��l�+��ۘͺ��7���$\R1��N�w8XѴ>���p�y"�Q����=� J��%9��)k����cJ����A�^8R*$W�����6��_%�I������$�{�j�Ũ���PVNZ�$�{�N�;�?<;fT�$i�hU��T��`�BUVX�T�I�����*V����O�;��������ߞ㚝��aO�L���-��`ǝJ�Z��z��{�RD���;��Tv���χ�N�Fe��U��u������C��*0mB5�,%G+|��?	f7��ɽe�BdaZ!ץKU�IЯ)O���g�a��T�f` ߊ"�>��%�>�|�a�*	O��V�1��ޜ�BxN^M_�/�{��dH؊�6I V�v�R���j������v�v
��{I�MOd�r.���:;��֑<-�%�0�4"�BZ��7�V�%�U����'�Npa,������J���O�� �&,���N�&PAp1=N�tڪ����P�U��|~�2�gf8>~�.�V|ЍiSy�^s:�ޢ���f@�~��4if�
X����r�y�P�w�B�%j)�¿�@d- l�$zhab�x����H����B�N��@�*O2O���y3���ׁ}7{�X����P�n>�%`�R�܈�f�bҿʺ�!W�8|����ǜB`�2�`M^���s�s�Xa04��#-�tgi=��4�ߢg����R2G<do��`��4J����c.z�g�-��r�r}�s;mn�,��=����Dk�n('P����q���+:�b�-�ͳG����]��S���,�@�����Dy�@����~a���S��6������H����z"�w��w\�c&*6x����I�]�FޑӪ�ğ`E
�I]��լ����?�X��t!��#��h��H.ᆳK%(g6wD��<�}lXT�����Q�aݔb�/�N	R�M� C�刘�H���iqQCL��
8�Pe���fF�P�aݪ!������95�U+!�t��U�L�p�n2}@[���Ȍ��d�rS?��B����Dr���I-�ջ`Yy��D4^��P@�YRg��d<y���b��>#�g�!NH�xی1��u����=N���:}�IFQ"�JVC0���ؑ?����5ϊ��sV)���뺮^��� :�H��)�n@{�u8�m�޻�*W1&���kcQ��J&|a�NT��5������W�2Z8旐$?(�����kI��i��-�D���46�v���:�N�hJ���(ht�ex��9�C*�Nh�e�^~�����9���F�&}�p��>��� ��'���^�*��z����wۉ�Uؼ�< 
(&�~K-�U!�=G:ğ���9:����ː�-�w�1�#�>4P2�e��|sҩ���jֹy�S�a��mp��R�te�6�3��.8?�C����RNT�Ix�kV��q��s7<��K��D�~T2�^��ҟ#NB�o��(0�7�V\�x�vQ����j.�yn���wgmh\�`m����Mu��A*u����7�2²���Dg>�����@�,9/�u3-�)�Ӵpj�rr����:���
�L���Y���7�����ꀨt���g'wcgAXڝ��6_YG��1�7\b%�8�dj'�_7��(�6�w��iX��,�U8�'��{i=���H�&�' w
H<r@����5L��F$9͋I+�J廟���cb�ۜ)G�ݽ������t"K��/Q�|�6BF�$6u�*f^�T07dY�?�v+s݈��D>���	�z��\1�����8�\鷃Y�:&�F����i�+�Q�Z���u�*�צ�*b���M��e\��g���?q� ^�}��z�������Z �ߜ����}0J))��vhv���M�s7�]ҍ���Zӗﯚp�ߵ�F��R��L�˧�W"�U�ʶ��=ď������4r%�t��t׶&���`}f�EYĿ;�t׶��������(���f�c]���l.b:���}�ZT��M!?Ï��?*83��t������n%gu6���&�l9����˹�"d��C_F���P!�T�A��N?	O�r�Nh<A��u���Xd�m�3\���XLI�4Y��w�#^M�o%f��ԉ�¬�~�g�+�0{��Js���Ϻu��?B7���B�n�fSֺ &o����T�&q�CE5*�s&'���*���y�'�-�N���.� .>-���=�W�0��:9�|�_�C��^���<d�y�T��j�<,�~T��]�Lb�v%��y;��-��R��M��|*\p��9~&�n{[G�� ���SSz��tv�0� ����VǕ����.|U1y`���f/)E���ڼ����l��u��0 �{��,R��Le�HG(�R]��U�����E�PoQ����Y&:�Z蕽\?����V�H_��"G�@�lU
���zE���V�E �,"U�a���O�Eu�@���IVCH���v᷷�sx�I;�)b�Z�䋮�/t^�+ɷ�﹞��,�\:I��	�?�4u#�q2�ڹ�Rr	Po�X�����ˡ�0>�R��c�Ǒ��V!d0w�5��Z5>��-��l�f����άF����|=f����~jP���2�L5�w�h�H�_.�T��B�^�T!R���5�G�Zv_#cL�ʎ�1H~�0m�����>��v�>vI~��}��H#E���������R����y��+�҄砡_)
��!�(�Cr��E$���q��fBs��u*�p��	 	VՍӿ��
9v<�)h���K�}���=��͒��6c��
jo�׭��F�OF�~�aτ�Z3 ��b�o�ܽ�_'�t�xK%��)ڧ�F������R�Mb�����a�,|GLm�pKw����O�� ��2I`�N�r�̢��2)������f8=?�e�	p��ԥ}Ѕ��z��m���o 1E��[���_����$&2�15�1�7T�͘�6Q3������i����k_�b����4��ڕR��[��˃B"����[J]�4-�Y~qMM��q8c��uP��0x���N���ڿ���p��ZD��FW����w��x�Kr%�c�k�yQ"3䳐�6�@<����N��Z�m�`�+s2�.����n#)��{!
���6��?
~��2�m�Z鰊њ��ۂR���̀�5�͔kd������{aV�����z�
\��%Yy<y@(�B4���Pw��ſ4`���n&#��NK�s6�{�VB{���@0��q�:}��+8�˄[P���*�ȣ�)�mteZ��i2X����![� ���H�yn�+��~ s��~����!�FA`$,������	��ѝ���ͻV:5�e�=�T&�D�K��EJ��]#����5/t(F4���֔��dk8	%Ȯ@��Wv��-��n���-��}��s�k��F����}W�z�8��j�'���+l;����#`F4[�aCv���U�ߡ���Z�8̿+��
τ����w����J*�٬MU�x
�_+��+����i;]2�ȗ;EZ*�O����fųTVv�b����٤ǜ~I{�̲�+�ds�n��s��볪��K<%���O�pR� f-)�$#��3�a��"����4(*l�M�)�wF���gw���ȩ-ل0�$�h�1.�B2&�7�x���r6���������r�ʲ,�ˣ�x:]\�)d)G�d>�W��������� 2�l�.��� ��e	��fv\p����S�=��<rl;@�aX		���١��sSmH?�����+pIr�v��yj�^}Y���〉��[(������l�ĭ���b�PH��=ص��u�Yp�^X�$2?פI���Q���B���_p�̓��5tn����I�_�+f@�U}3ό�<X�vX��j�~g�	�@�Z�B� �O*n{��Q��;.���;���xM���3@�8��^��"Q�꺖���|-���?�a�֊%�Cd���G�e�.R&�b��E�͡��ɒ8W��.G5Z?;�5�����ʞ�w0�{�T��Ȫ%k�TDM$+u�S��#;����®�WUy�n��g����c[�]x ��%���~ĕ`v����Z�L�e�Nӏ���ކ%M�����ԧJd�N_Y��y��<���.��|v���&F�ͻ����6���H��i�/��MF����<��䳬(g�&ë�*��>����R&tZ����	�]�~���7C�NH��J7K
��E��:��H�o�;Ux�CM�&Y�A��κ��F�6�Ѫ>����;Ԯ���̱��+a1%1��L0[�;:A,���H,�ay��h�@Ss�y�lꍓ�5��G��K,WS�ߘ{ zN��d��Z��ڔ���~�Z<KL�+�
�i��t��d
����/���{"jrIR� ���S���`��f�A�������GyX�V����e��`����K�[Q��Ć�Qu�-_�R��f�pr+Owz��k��[���kz��*2
�V@!�t�������e,/W (��+rn
�e�Hg)� 4�����v�(1�a	F5�7�q8@Zc}�;���������،!��,L�dD�TG���.E��/l���b��I�L��.6����1�$S+�8EN���,}�(~���TSl���"��Χ4SP9k�|��Xo���G˙��4�VA�����US_,����y~(�пiRtI,Éd-V�TS�7#2��I�� 	W�	���2u8�]�� �ɣ�h�t벽��|g7*�b�(�M
�l�I�R� ����n�AE�CP�tֵif���&�5-8�꟦
;=$�a�Y>�[R�~Ƃy��0Q�i��<�`�]dO'�ၪ�n��^%�ݒ�n�~>0l+X~��K�r��� /B�gي�Q�(�a`�\�ޒI�����F̷Z}��C�Ѡ�J�6�xP�}��^nCG�,{U��l���2i�e{�a*���rw�DH�x|_��5�[9�U�R	��������	&N��\�|�q�[o0��0tǓ`5�)|��:&�g 9�ߠ���.cw�x��f�9F|��/�>��q,�f뫍mד��P��Ǟ7y�8mm��p��1�W���
 G�F)�Ǩ�|Ci�zˁ�
,�����N;�+а&�7w�"嘃��VRs緵��0�ߖ5s�5=���5Y�&�3�wX���qC��,N.���R*w�nx�nA���-�=��a��_�*P�j��㷌kPd������
�vB���D�I7{J_3�Bq#�8nL��� $/r�=M�.����D�m?��(mp�ҽ@V����̠�栏I$#�d᷆~E�M�k2x� Jr~C�*� b�wˤ�jF�|�4z�K�6�T��տ���<%�o��&:�vˉ��}�v�vY3��c?�밢�ń�ȼhk�C�WgB��LgE"�Z�Tp�=
��ѩ���Gb�WR�`1M�4+���F��M��0,-���xQ?�R�k��o	�7'aA�гa����g�S}>�Hю��B�b�G�⧙�$A�GPC�v%����g:]
}��
q�� uAJb��2��=v%:ќW�Bb�l�:�|��ڵ�FJ����"�*��+~���0���� ��K-�{߬ʞ�%�%|�r��2T��ˏ�9�p�_
��Q���+��2�޲��t0�����"�@J���|.�����K<�����~��	.?���:GzSy�ݻ�籞YVaT $�}���6��`T�SM�LڈF�3@#@8"O�<?S0=�%H1*�T����3,ը�#�����Ѣ9g��
��C���dW�Q*j��1���q�d�#��{�~4@���_�Ø߲�9�lu%��`~V�?����#Bgn~�8���N$��U�>��[�s���k�e{�q�T�3dɂ%�ʷ~����,ɖ�M��r�J�����>y�O�lZ��8m�5�#��0V:�d��$n���$�ƹ�f#[�MիGڂ?lg:E�,����Y��k���PBfY�tQ�J�l*S��P/n����,ʮ�O��Z�s�dM7N���\��#��-�5{Ќ��p��9�h��\�[��mԄ��b�|���9]'�V�0���z� ~��r{�-��*�m��FØ+��>�U�;F�L��|8�-��ড়RE^�������U��|w�X/|R�
 ʇt85�C�@C4=uZ�V��\9�̠e��D�Cx�{��?�D��d��,���Ĺ�&���	-pO���P��� pE�p��0��Y���O1>���Ȣ��Ŗ��.���}d��Ŧ���Ή�	��8��w�~y����m���g=7�脊�3�8Y��,S�$�2 1z�B�����U�5��J	Lr_<`l�e�u;�"T�O��N�.�� ���7���[�>���M�����L�o�����3�Dq�lK�>��wxo����	��O-�ǇN��1iH���h�lT^OsDG�f6��̭&��ja��{|��z�[�.nn���c��r�O��[�Ⱥ �@�EJ?���'��~���Ɍ�Z;R�J��.�[!�$�b	���9��O�;r�� }|0��^�'O,�7���{Y��H�C��_�d��R���
ƙ��JG�'%�[��9�_��2��u��d��9ߌ����l�R�
�+̼0�طkR�9����>LϤchġ���(BW�.������]���fL���HO�k��shYb8qhE���L��g7{G�.��VU�j^Ci�y�Rq�0�Tz��E�F
�b&��ո�gK���]ZZ铡�wLW����-(�Yɛ���oŘ��]I�R��U��qp��Bn�X��Kd���~9a�̝h����)D�cp�����
]����V;�\������ƸڮFȜy���-V��،�3(h����� �߉AÒ�'I��(��7U���sD��'!���3S&�c�,�l�?���b�_�U^�F(���xW���k5�j�Vu)�,��eP(�����U��4�;=�A�~q&��_��i�~3C��5�dE�Ou#�T1�GZc,u\3�9��ae�	�x�z=���ӌ��K$�g]{Y{#̪�e8�u'�bJ7-���H�97a��d���}��!�A
mV�,���_-�D����>�_�y�8W�3��Y���ע4֣��_����Iq;-��J���ͥ�b,  ��bkW��#��z��o�����^'�������`��Pg���d�W�pINy�ΘhQ*���ѽ�o!��>��!f E��\�;�r8J��H�y.*k�@��������R��^�]j��e},З�� �2|�|���*Ɖ\n
� ��m=�7�v }�Up;W��	���Պ"�I�bRU���
�F�|S��n2W��x=ӽ�J*s���кU�`,��KYlW��.-�����d��)�ic*�&��Ը�In�.Z��F�:/{�e����JdA��!����>����A�+�e�bN�3s��m�,��[�&���R	�d3��rӘ�=�T��u�����;�b�XIg���B��mo�� ��	�!����e웯Ge��oĳG7���m\��0���
q������:Q�9���oR-g�jd�ۑ�dY���%�3@{ۊ�`�=�+wn��|^����M���h*�1�����r�vsg�1�.���Z]RN���헛��>kH����r�c_޾(diв��\މMR/Y�#�r���kM{9 4�K��J�F^GԔ#0j�=�ˎ��a}6̭�9�݆�h��,��]�g����z��<�N�s�ۘ��Yf�)���Ē!y����mB�2��Q��7w!�.�a��g�+H�D!#
�����~�!��j�Y�ʨZtV�pբ�:��������p/�k0��9�LRB%��gz�і��F���)��A@8�m˚>R��z�d�{p��$�Π5E�C�Р�Y��Ț��8�qC/M�h8Yl7'ӜG��u^~+��v��"=��ڸ~8�����~���ca�/Z��B�5�-�l�h��$5q�m�*�ݘ��`���%�U���`;"�QWq{��ޘ׵�^C���	��aU�:
QI�wr;��|u�N���#�a���AY�
�mt��yq�$N����"s��L��2la��3��x�cj-�	Uh��81ɭ1�h��&�-�6�И�O�'ƚ\~+�r�&G��k����cA�K�� !W�bƬD��"8}�P�<cdM����E�g9h��ɑ�%�y���!���iLj�/}��̄�%(�^��_E����-ş�u��T����E��zLJ��7�c�t�;#��H*�teMRah�����ݿ�q����R��c�!�����k�@���|�2l,�̠��&�.  �Ց�r&�$�9��ƛi�U$�]�޼>�J��&��Qw��YR��"F�>/��]�D�>�aÖj�j�E��C��VËF�C�<��
���@����THc��/�YF�ǯʥR���.1-	�sQ�����Y��)���K��|lUf%�x��Q�)A�����׾G��!�I�:�?�,��.��H�n�Ķ����9؏�a�ݞ^&��׌?P7Vӽׁx����_���[ؾ�3���I&��0�;�,���ω�5�[߲��^V�O�����ٮ�?L=��%�8ϓd����R���3�˲�5÷0�54 ��	T�C�z��I�Z�9d?EW�W��]sa��RԳ��<Ieyʞ@��Ē�;��������W��rvt�#|k��	B�:l�ʱ��w���&���HB �Bo�[�1�*������Հ�����S����T��y�d���$E�q tbu߿�� ,��>�\�	"$����Z�'ڵb���P��/��!�I�i�v-	Z����f�P��=������I��~9��0i����EY�@����1`��8:-�?��r�n��
;���&��e�JK��ޙh�������0�`UD�z^�7�����z'��/�7�߭�/���7�W"D�B�6�� 9� �^��)^0G��})	?�pP)��Yi�����|:�LoU�aM�Ho1��`�Pw|4�Ћ�>�8����
��CՠF2�y߫}�FER!����T𖅵��7�iK<e6!3�'�{��lTz"Z�2�O�)�x���K��tn��hp(����9����6i�����h48@�v�CF�:<gfO�v�� ������qe9����1�[��?�V�<h��)��<�`ց	ϵk�ܘ�*����r:>/�盟�{��]ƙ +��M?)�Rq'-��ݸ���T	L5{6
��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� �����ޜ<(��l���R�l�iD�}�ŭ�L����6���8ﰘ~�Y�xI�h
�]�깵.�0i[�!:�N��~#<��3���~T���Ođ[/���e�fҾ����_6���*��"�������,TD�N�O'N��q��)����Q,�剺h�L�7R�*g�t�;�nG8T�����±m��d���}��٭;Z�����2���_���w��q��2�=��|׊U%|ggT��+� (`@ZĹ�KؚU�-)��w�)��,�g�A?�1�}��
̠��d�9���`ힸn%��Qq�a|S$���Z���	T�+���v?u&Q��xO3NXz�i�A��3A5o��k[U��jڊH w\�'�3�e�!�����(y�<�p�3N�.���ɴ����2_�c�H���[��#&n�D^�����E���&�$���5�7J��,��W�yk��p�}�/�9��z��l��}���S�����Gqz��ֺ� �쯺���h��^��SIm~ �����!V8=8�&1.�hn���Γ�-YК:�i�2�p	 �&7�ONz�M�?�ѕcДe��A���4�"�f�o�kG�~z��B���t�mU�.�u��j�wy�ѐ��eЧ�%\�Sg}��|��ѕ;)T`�������-��$��b����w�M����]��M�"��Ɣ�B!kuy��*T�Y*]�h������|�W-b}�kH��tw��y#�N��{A	�w	F���/���(ݘ	[�"�2�|\�؆��|	I���!V#�7ȉ�%^�j�l9%^�sw
��y�׍���j���d~��L�"$FB��t�G����G'f=-�����a߼�&��2R /j����B������I;.�<������Pk����5�&ɯ^�Gv�Cѥc��:+�
~л�ㅮ�8����.I������Q�z�=!�ۖ�~�E�Q]][79�r�{f�û�=���J�^��"Z�BJ�N^1���Q�h`�b<��JxGe޶��Py��h�5B!�/�,��׳juf���d^�kmZ[,͟ߊM�e�r���ߔ'P�M���ov�]��4yj8(����	Yh�
/�/Oks�KX��oan�����x$�h�h5��R\�/��*;�A Vs:굻l���֌���g���y�Ȱ����߂��z��{R	���~�� �_k�d鶔7�!x��d�&,�y-�Ѡ1����A*1Խ ���s�!K�� ���T�)�����>��J��F+����7h�rSb���FnP��
ÜO�O��0��H�AZi�,����W�<e0kz�vG�j�B��S���RR��v��5�c�w
7 ��)���V�9��@<ؾп�9S��ŵ�^�;���OFZ*�E���Dz�=Y��$��y ���H�n�?/�Ķ��ʙ�W��<>m���'�u"$;�,<���:���3�m�]�YU-�":6�1���}�x���(հ"X8�;�(
V3-�~�_�Wf�K�U��}�[#B(|��=�w��8&y��n�Y�:���Q��$��Tͨ��kJ��;��M�\mJ�^⯬�Q��b�7�[!�����u�s��v�pg�]���uL&�"Nч�^�3�DR���ʋ�3��Y�8�Gw5O7=�u�o��5gϦ�ſ�>M������&�v9
/@�.v������,0��-_?9������%(�J�ל��zN���	C';���κ����� �X�5f@�\5�V: b)2�~��kj��eO���f���a� k�gǐ�,LLxdv�$bV�V��������N�������B��v@�noJ ����`S�������τF��Ǫ��XZNr�ʮ��Gs���%/8��B[��#yzg���B����@Q��9�a��s�S��a>%��~�<�+��n~0�֎@��-x�ɲV�C�x0���z|�(��a��_xhAI��5OU��m���_�������E��*��z���&U�6P{�zy�I�C~Ll�F��]w����ª��p3E�SДV�
2�x7lS�4����{(�=���Ty����ż=:�S%�����570r�q��Psn��&Eu��\�گ�{凼�.�xY����qP����o��N1U���Rf��x���G_햐�qU��9�QgR�����wԉ��%�x�s9����/�+
.g`�?@"n�ZӱJ0�x���zl7#:KH�y�<ХU7t�bʁ,��|�)�n����0Od�ܮGi�|��U�O��+-�뤻\[%�&�vi��XCƩm^������`E�·z���#<�	��Z9��恼�W�bm}���a)���Ǟf(��Ӛޞ�d��p�z�_�F��I.�-��m�<횰s�ZZ����"օ��t6v��rn+Y{�S��Sh��U��)���C�Eb�;�Ҙێ��W	��:)��+u��/:������{��5��19�)�m���t����S-)#
�mq�[x��6�B�жX]��t�A ���HJ�HS{��E򉴦J$@�iR�^O� =�#BcYTWϙL��
�'�쓷�|k9"L�����x(Eޡ6Ygd�t�Y�6X���>:���+/��!��6�>)��j�e\8�R��"��O���ilAe�4��:L7���f�vICH|�9�5��i�K=�tӽ��Mu�f[�V�1X�&�p�j��^W���_�r���`�pP�D+�����I�ڑ�3�&���z����>`�"�>��Z�)?�:�%��Ch�-r�򽭿�;�b$6�)��ȯ*L�_~���x��`��4��q6�K��;3�{�Έ�em*qX5�e�-ۚN�kg��t(�������Q(�����>�M��d�p�޻�tV:�k��S���Ln����dP��Ud9������{�̖��=����RhM%/@U!`>�t�V�A`�k[AS� �!e?g��2O�"�oH6=���~a�M�s�S�`�Σ2�V:�]���3/�����{�^���0~����Ph�1��eL�)�I�+d���m�tA�
�oO��.������6��q��|�Rr�Sx2���Jⲉ����5�ݻ��{� be��z�M`h5,Rnnfɻ��}�^Q!A� �SU��zY��qt�, �y��8���c�T["�Խ�$8ܼ|8�`ј	�S;%��%�#]5����,EZ��'8z���h�h�AoE(3��]KLO��0tb9#f�Ec_�p���&���k*�aꟳ#��:}qne^�	W��t�Ӯ��(���E�jL�JE���ҷ����Q���1�9a������y�>��}��Kf�	y�-{8_7n�>Ra+%雈Oy�n�B)!���C�Oĕ�c��cH�]�	]ǿ��!6a�m�dx���qp�ߧ{|;��V�mJ<T��q��u �K��頎`b4ݤ�B��vZ{����=8���}}��$������=��p{�0�E?A}��p�2�V�3���M:��9��i�Ehψ�}�alO�o���"���!c�a<0=!X����^��@�Ӭ��Ճ�f[3C��>(n�=PXG?��	Y
�q�����R��f�8HgZI��h��@W
/o���CT{���;�m�$�����)� R�~r7�2���3��2��_=|�@L�r�3d
���A8����:�Gd� &�SfCRJ�ґ�EC2� �0�2��ļ�R/A���q���S�'#���-���PV2��l��u�~4<a����(�U�S��;�ğ����8�`�濮��OM��6?�xR���?��wf�@�q�	�z�7̵2,�U����f���ʼ�#;?�n��+z�o����~�"i������ �-x��hC��"���`��ޫ�6'�Ý�g}Ƶ|ka:����*5�mJi�j�-�D�,�a0*�d�f�;��ύhCj��.���m��DX�Hϲ��Y_]!��Na��� *�SF�D&)I@l-�$��zj���~����k��K>S�0���M/7���8~ps��&d'h�sR+�<Q�"�`85_U֚2�6�~T��!��U��h��N ��-�#���$s6��P��wHbs1 �6ͥ/��R��u3�Hf���2O}S��/Xk����>l�VU;�{x{O�!�8�خkcʍֺ�
���VUУ�$N�V�����{�DӆM f�D?w���̄��\ќ�^�����F�;���i�J=�Q��";�6��3}y츴�O���ކL#�f;�#���ܼ��R\t���8��F@�J��f��0˺q�G����b��
=��N�R�Æʳ��u9��{�=��\�BE��bH�[���F.r�C>:�迨ռ�������ǹ�:<�јB�� ����[���:)DD�v��X����W.r�J�IDao�|W�fĞ�U$�:;	^��j�U����[���]��9���t��r�o�m��	���F~�O��zo#;���C5C��N����Y�(���f�^�u��x)�S/�$3')�f� +��o>fҘ���h�C����]"b~���s�^yd�9�O�e42��[	D]:��t��(�M#��\�[�̐:Zph�u��=uT��UƠ ���ǵ��� �'{��R�[�_�R�I@u'~�,��;R0���99|5*M�i�S�ዊ�'3�J��
�|���3/��a����޺�۳m/T�2kE%6���k�Z�3�)B5���r�]�**��-��<H�`C�v�Y`�6�h۔��a�l@{�`A�����ӡ1�Ck�9����Y��G� b�;��ɕ�����mQ��L��3�V���c�����T���~i$3"��;��tD� �V*���ZPhU3���Z� zh�-�/��Dro�\M+���iuo�D�������e�͆OF�2Ɣ�|O��e���UֆtD�1�&x�+:��#3h�	����S$�pP�"�v�nY�9�>Q�IὯz��,Z
#֯
� =��GUUe�I~�	ް�-�)��q�&�н������Q�������B ���A���>0�C�� �����Z�v�-�m/Z	���_�.i�i>\7���I:�ph;v��ռ)+k�wa<z����@�@��/`�./?R����yن�F)�`��xHepr��ћ�.r��>��G��D2��C�"(ݐ��>A',��s��z���;��;���R���M.GP�����BZU�}���������������w�.JB/=�lϣ��(��:��z��-6h�B)�����̃Mf�4�4l��x�>z/e<��BL�%)r���Ú�Sz�{�uI�&�$����ŬN�~ǛZ�=l��9��̎X#���P.����у(�֠�ǹ��,�h�5��L5(~kg�/Qs0�'�m��{U�&�Ɲ��nN��I�B�.�[--G����[��G�nI��j�=t�
G6z+[54��G��.##f�k�����C�v��w�k�F͡ZxZ��?�bdyQ���[-��\-��J������V>��v�c�m/O�������	1�ɴ]���3D��g��r[�wm��?�i;
�Z|��2Gm���-��>����_��|�Ω�̍��-{7nt���qrX2~A��mPʭ*@�n�M���M����-���A7��IF�~��G:����m�۪	t��:G�CJ���tm�᯿�I�dt���n�"tl|L�)��>���&���m5�^/>�GzO�ݘa���k�ds#j�+�rI��E���1ԃLD���K)_s�5�4 cG$\[i��X����\�=��}��0Sj4��jyV>3m����M�������2�.�۱�Ж'#�h���m�e&V�i���Tu�p�z4����SM�+�7��š*)Ǐ�z��p�4nf��%0�ϩsN�#gH��J�ÿj��Ǵ#���;A)����"���9�\��ׯ��io ����K�)�w@�I������k���������Fn�k�+@�񂯉l�OǕ�Q+���L�� �5����6�.ˉ,���K����hu����ÞIc՗���W��-Ag��"sg��Q�����嗓�'տ�W��@ct��\��9�<��UE��	K[ms���C��R��I�{��c0�p�qNk�<��{��Xmd)����L��>�X�S$�����>� �O���O�����g��sh�P�Xb���NiԵ��;��4{�>���ucyg��y����ΖZLm{�L��AsR�Pظ��NC+�Gs���,��&jg�'�W�j�TY��Z5��Ӆg� ��Y
���r@Џ�e�h��1_Ϸ(=f�PV��~�+�u�f�ٛm[�zW��ϲw�J�D��0�'
�K�i��
���/yw���J���B�Q@� ٕ��q�����h��*E5I�0���YW.��I���1�o���^��y��w� Q��
h�p�ב�����v�"0����2;���#Kp�H@�;�Me����iF���𥫣
H!顸;��{G0��4�_|�!��sᰑ�lL'�ky&skg@ݔo�24��z&��rɤ�T��6:f��Y�	[�A3��}�ꪚ0�U�1����W@���1͋�⺳�-:�j�+\O�Lc�͵R�ѓ���Wa'Ϳ3�٤2F���M�EJ�s���+��-7�/����j��A���X��J�+�vO�(���㜀�,��a�)q��e(*-#�p	G�N?�N�,8f�J�  �L�+I�^��X~
�	�#�Mh7��<~�,N$,Ҟf�@*)�1��(|ȝ!8_�X�pZl�n������a�� Q%fj p�%<�]c2�3�VF�##�h}��Ρ"g#��V�J�|a��%'Q��,��J'����Ĩʖ��!�d�����-��f-(~(.�e�W7���y+�!d���"�2C���Zʵ2�r��9V%E��MMk; �tKx���U�.�e��4��~�d�M�a/BZY^�QqZ�+�����i6E���8���m��U�աqb��1�P~� Ē�J�Y���G$s����#���ۖ�g�\+#���az un�s� k.��Ai�/�q���N��v��C^>��w�^� ��G(9��b�ڎ �O��Y��m��B�c*�0d����k�K��ݮ5���o)�p�(��W�1�yxܾ�-_ل���H�	���lZ����;�8ZL���x���Σ�CR�L���U<�ڐW��iC��YjF�ʤ#-4Q���//�e� Q:]���SL�I�����!�
�Ü�7�!��X�W�	M%�hWY.Nc�D�P����~MP'�>AM�%�+.M1�U�/BQI'ޚ��:���OՓ��u�/w��x��XkD#�`���M�y[���2�� �:�.��TH@,��#5)�� ���N� �A>�o�u��v̠k����H��N��!*���7����S+����㮭�i|�~DQ?�ښ|�b���I�%�~��ˍ����\���E��`��(���5�Bk�0C0�\SOlt�s-.��K��Y�׃�����XY0�ڔ�I�q
��|�]�*������VoR��M�4��H����o�;ӦkF�隇|\��EQ����%x��k ��yVCl�O(�h��@���_#6_��y�7��'1��Y���h(f�e]y���/�ӟ�q��,^F'��u޾�N+|Α+{����w��ydl���d���<ufyU�#�� {7��(3��V��87s����3�M���0�q=���T�?�{6*�v#s-�r�������ɏ���RG�n�Q�A�� ^ӽm���̸�XZӏ� ��^��U�@o&�k[�}��^{r�9~�����V���~t�ILU��%�j�5re���]�S�%�K}�L���y�+�w�
&0��f�$m���IE���Hs ����o�S��>�?H4LX�T,PB�;���<��T t�c,S<�
��z!1R��鮨�abjcmRj���d�0�K��I@�[�9��N�]��X���u����zz~��r
A�f��~�tP�~�W��\��j��K�ٵs�m��z_Qlr���zµ�Y쾅�� ��Y&/�-`3�t�WڴnϞë�| -dH�f��繶y<�P;0�U���YU`{���P"�3���O�4���M��[!���8ۜ���C�"z��f��+�TЅ��o�$䈼}�Qy�2��:��g�-/�����{"�y�aT�Ͼ__hwd��Kz	w�M���L�R�֍,|����K��}�����L4��*�/O���fOL8���k�<�U�/�85~�L�{��qGWĦ/Q�,>-33��tx(��?Xܯ�����{o�D�iy�ހz�o���	����#�����p@Y�޴�I�1��^y���	���~�\�LϼE��<J�u�����csb����Z3�a�������>���[���3S%D���?�j�k��N��w+[�x2����¯�e���R�=��DW*�%� \�ϡ�m�x�6�	sH@����)��zP��iD��a�p4�κ�+�I����=���JTxUm:�g>�kZU0f��urx�@�>�)$��|	$v�5�+{��R%y_8�v��j@��������CMq�h�;�tf�4 
{�k����-����7�Oث�L��h��~��:��
>h )Ι�y���T*��u5����s0�K�eR��� 3F%�5��@�y�<�/0�K�ТP��ωو�KK���'�S!d�j̏k�ns�2bI���1�#��2���!Hc�=^�v<�O+��;��4���<^ox�ǰe�O��D�ϿT�����]S�@�#o� 4.PD����	�.����]G^F�g�v����&���?���'���$�O�PG�qCR��x���7I���B��������BA7H�*Uϩj*��%��c�W�?��n�EpmѦ�U�Ǘ��`㗷�ލ�vҊ�6�^?Մg�*�ӹ��P�QO)�X�J���I�@-��Kꢛ?֐��t��{��I�b�h��A�ǡq/�F:�C$=9 ���^#�p(���U2�u=�l���'=���M�&�;e�9� �� ��Y>u�)aS���xb��n���a��=W�����ǎ���_�Z\m��T0`*�P ���8�TY��@>��8�����	��ԜI�$qQ��.E�z�2�0/���w-�nG�����}&Dfݢq{��I��ۑ<�~��j��5&�@~�1��i>%uAZr�0q���p�VX��\�F�L�\�� �P�bR����1 @ȣګ�G�UF&���'�|f��������t�y�{��Z&{�Ő��6��)K�xw����!��d
��C%�v]ȼ���4a6��yKEE�`L�D���|��|���G��.RF���Of�2�.�j���g��ؗp�K������p��x�e�c�͎-�|�ž��%e�'UƩz�+�q6��H';Ijk��vÕ�n�o�u+
6>H�?�.
�"Ih�G���*sBJ�g==�l�J{�8ѵ���H���Ĭ���yc���x{R��<�7ΫK@����W��):�5��!]�a�g7��f�p`5;�U�z:#�2�;�������ǈ$��DnfR)�ƴt7����aWzLK!|@C�"M��ΣI�a	x��X�Ǘ5ER�R �UJz	�G@���_�XNa�<i�^7�ˑ�2����P�]'R�6���j���s�����U���wSS������a�Ϝ�]/f�k���!��=���o�ڦ=^�W��0��� ���A(?��vdξӎ�H�	�xbN`s=�s����Q0�>7�	L��+���Sj2\��$7edl_��s�ܙ�h#����r8���2w�|����kYf�����0���� ��0̅sW��Þ̜�.����I�8�Z�Y�,�rf���8�4z�uu��Gy�_*�QvN�g!r�o�"܊��^�-�!_��;�p� 6.<c1Y�չ�z�gB�~Ļ�@�±�bdv|���"����n묵��.}�&sB޽��O��wG7]o���D|���>�c2�,KR�E���`��C�I����נ�%:�A�X��� �ڌ=�%"�R'���2_� ��ڥr�Qf�7����^O�<{���"Iކ{��BK�Z<ϒ�������!z&�_�|V5�+ypY�J��-Ф}θ���T�
9��$$��_8m�����G���J/#�T&��"� }��͸::�����)�R�4�����ƀ
ψ��X9k,�E߆��
���C�]*C��$�]�s�NhlZˣ����]hK�<;�z�~17+�Ham�ȑ�2@�7ٓ/�u ����	/w�Q�a�V��W\�W��?��/`�8"H�g�ѫ�`	�n������M{	�_�����}�_?n�u/O��F�3���!̪�ߢ1�.��bA"'�:�k�L�HQy�&܏��ΩXq�V�	����䏧j1��c�ݤU,��B+H�dl�4Aӥ����!2�a�<Hd�3=(�n�}ęo��]�%������@9��/����K���i '��4Sa�����(Z�t��f�ck�:�
��
[��̨ȍ�sֈ:OW�)>+V��S������Z���c��M����4c����b*r��h�KZn��{��)��}����9*�)f
�M)�>�D��>TRVm���kjD^\z]���L>�=6zvMC�ik :������N����1�B��*w�z�z���`�m���v癮.�}B%N�j-e�5D�=�\'���g��?�{�b[��\��g􋕨>j3p�w�>�i��jew
kE��N��QU}�f�C�I���N�x�:��`�am�{��=3J��,i����ݼ�b���X��f��Z?�s7BO���L��w�;�hn�
�iҀs�"[L)���O�}T�Ʋf��ܱs2�&��yȌ�60�����F�9bx��r�vp,����Ug� �C8n�U�(�>ќ4���u����g����Q��kv=z8��xl���J��y�b+�?z3�$ö�WHe���?@�$EQC��$�$��<&(�=����2�&c׈�����;ݼ}P�^�Jf(�8i��
���&�������]��=q�%�m?�d;y:&Գ���F��6<;��,�(;��1��N�X���و%�%0`��TsqX��	�C��6�1����FM�ck�"�b����>���U�ۼ����-��2�_�X��6e�=�F/jXs��9Ә'��B���g�?���L��,$0���:"�v�=�͕r�j�	�T��a�a����|�[�)�/�Ʈ�48��S���5n���C�{/��k��6�m1�̈�� :e�w[r�%�! ��(���H]�+~�q��\v���>m#���?Ӊ��ȇm*�6A?1ބB]A�t���N)��^W��wpM2o y�v��ʍ��K�$R���(OJ}L�A�G�U,ڙ&x1�8$���Y�ۂ�_~M��]q+/��y���۟��"p�>̺�J��I��u��O:���`��2M�P,y!kP�=oݙ�A¡���@��Y�^!����g���S��哵�h@�IXB
���?���&0��'z�;�,�Mu����7/ẍ́z��;9�~2����pz1���O�f�h���HԮgL]L�P�SV�.�A�!�b���EH[���o��w4����Z[�&D[v�fC���|.�NU�HZ�ిv�il���)ܝ�*�0�}edn��|�P�n���'���Kǆ��X QY�ƻ�!
FM�1D��-N�t.�esƪu
�J� P����c�.�5�]_M-!!�D�1o�}u��f�*'�F�-�Ҥt�%)W/��f~ѕI�j�5GB����2l�)��f&I ��{hKCP�q�N(��k�aL�e�����Po��:�dl�G`����D0�K�-����,�\��X�/���-�_���ޣ�����q]�!��+
�,hr��ѱ^_�Y1Z3jāU)���0��*bt?��_P��L��i@S��?�-w!�eN�8D��,�]�W�i���Z#��&�}�%���/"�s�@Z�&φ����	��=�b�VY1����u���Q���T�L�S}`�erx�b#7������P��lZ�EZ0�d釲�JXU}�@S0zh���bK�~b*3�HS܀�:���9>_��Q�!@D.�jūF�5���8�	|@�jv�9�"�].�UC�!�y��,���q;�?�^bjQI�t����庱�'ڇ�An�����j��F���C�+�U=s0c��I$�����i>��)W&E�y�����ӝz���N��S�'L_��7pP1u�͐�w�C쒘����F@�:Gnp����*gP"ĸ�d���|*Ɗ�D�������Dݖ�M��N �B��ô�S
`'�ZL�K���雿=��m��'���qTx[
JXv��O�B-J=�7��E����*s����v�kn�4��C����=1�!��Wޑ��t��Cz�E��3�v52�D���+�W��S̈�շ����%���T�j�p�A���M�0eQ�1]$����� $�  ���N={�n�x_< �r��ٚ�ʣ����ȍ�p��}�ܽ6���&K��)�ٹd�@7�P[řb��~�����td3Ǐl0C�g�.��L6�z���HWs3_�N���\�9HGl384��c�'%��Kg6�����a���=�t��d�_,Q����nly�����ݻߪ!Qt
o�E�{S9T��" �������"���K<X|�����G�x�
�#J��̱?�,ir��'��#�˦x�v!�z~�f?bP/�0"�\���;�����퇋��G0*�k��b챈�龆p���l�[�`���;�Ж<�!{�n��q�����K�pr��E�"��&aҒ�T��k�Q��7X��Q�MsVC�Ml�}%����I�F$H��7B��B�Z�Q����~d'��7M��� �«)PߕX��F�N����pK�H;��̨��"��Pa[�6��C`dO��p���h>tY�EH���O� ���@�6�t���ɛ?8=�w�pċ��!]�ж#�W�a}���L���_���Yz��	)t�ۊ1�Ɏ���/[�H�h}D1@9�FP�ʇ(�].��sh7 ]�ը�,E̂�Y׷9�����|�$Z��ȠO��ks�}]��jݢ�x$��-�79ר�2Zk�u���)��S�"����F��E�w�(s�wʫ�;�՝Ia6���u� v�r[R�� *��ѰȽ�p�&�����{K5b���pwo	8�m�͞UR8��ӿo3�!�ߞ��"�~���а�65��y�sǽ\�C��a�X}C��K�:9�;��k��t>���l ���&�j�Ļ��J���Lz�_�8]�L�<��p�*�C��p�T>���y1�20�20nk�֕��]v�\���m�tx�Jz� R��|�jۚ4��j"��WS�|@��{r�q���� >L%�\�� �@�U�*��.� ��I�QI-�])~��c@֐��O�/�Gn�j�ܦ7�v.�X�jd]"r�ΜP��דF ����A��H�'U��D�W�P�n6k���d����4TImf�G����ox��ЪYI�#&�l�¡"8a�������q����1��wR���F��}⣮n(�E�J*�3O�T��S�k"����_�8��kY����:w`�(#Y�YmӃ�k�Bj`�^5~_�q��^�s��s�p~�Ay9�����=d�Ir�V>�},;G�Q��?pZ�0A��V�I`���%ޓ��x~�`�(�e�>j%[��7|����\�s;
��5]�P�?<ތ#�������r��k��L;�S���W�]Bs���AOM�.����3M��hp�� �������y��`�X����[��� ���������~(<Ç,}-�����.�N�����Pչ�ዘ�(G���P2pv�:7n!�w���X�a,�e����l<�����n���D`.%��my	(��!�z��!���!���ہU�a
^�C`C63Vm2)��dM���E0�����2�o�$�L��L`'0|�9>9��_�K�j	�[~O�Rϓ��D���q��R F|Z"w�h�Zu!��G�V�rvZ�����DTK� ظn$d�����V�L����#�B��[��B,*����[���X�E;�\��x�_ʣ��(����sk�l���+Ub�w��~�LIu�M�T[�\��L����M=�ê�BF�&�����S�+��j�Ɔ����F�����g���� i�C�^W-������r��=q&�;hGD)Y�?9��\��Y����-���#1x��cm@��v�X�*�vq��K�q��GǺm �8�P[�C�W��y�y���p��ݷ)IN��i>�|����!@���GZ���0H����v�-���^�ҏ��/�$Kf���
��J��
a�6�=_N=�U?�ֱ��@�z�"�j�,�������f�ר��ۅ��O�rD��֦*/&5L���<v��ꭝp��q`����1�a��͍U�� %�H��)�@]��탚�ؑJVb�,0��][�:����6*_��F�8Ri�T��Z��lB�D��9��%[U��>w�X�8�!G�5��@�J�B"���Ū�+��9�|0u�E�ݩԗ��J��K�f��D��#�Yc�/{_~L1�^�x��	�6��T��%�+���+�hme*9r��!d\�bC�v��E���n;�l"ù 7�`�d� ��'�
Byʀ��& ��E�i<�kJ�"a�1�M%V@8D���$�>�|"�[h9 6�x�}����^8��y�������N�ﷳ�J�d�7cQ�ζ�ǝ�����!צ�K��R�� ��F�Qf����Y�$v�o��c�C*��u����S�����@M@b��ιi
��hz�-�VK�B�Y>4�g�r�63�:�����m7C���T	�8����q�<�u'QM���yѴ�P�����i.���UN@ҽ�F3��?2���'G	���w��F�)�-�Z����ס̰r!��6�5�w��OB�q�PX�p����x���(�5��]�Yd�u@u�:rV���`ʺ�y'�*�qd�'�U�0`NF��n���'��x�G����6�N+��� �{@m�)�c ��X����"��N����r���*�nv�c�wY�/h!V\'���W#;#�ƪ�����������ġ�cc9[߫��%����l#3nF�9������20��o�*��K��y�4BߺmC�!��2��֛������0�a#���B�<Q,6؁���_@��ȿ�ҁ��_���b�W�D]V�ӟp	^�G�o�P �j�o�&�ퟴ�hĹFQ�?*x��A������t���mi
�4�Ad�mEj���A���Q9+s�i�9�B�& ^�b��PͶ��b��E���s�A�#�� �Ӧ��V$�*�x��D�
�e*�+O����;j�uJ�tS��Z�'dL�H��EMg9y5�Zc3��dz������v���G�E���ȾF�O���,���0��h{���TM�5FT�c�)<�+Y�o��sd�-"�J��D���<+�&������gv�p�!���9*��	�U�=����0JŷJ���;��B��4���K��Kc�����5蚆S0W<H̯uC[d��61�(��Ɲ� �%�^���*-�v�W�rI^^rYp*��{�7 &�A�y1Ժ�s�O�g����L�&}~���i<��$/�� ����/}��Ȗ��m[k����TMI
ahL"��C�����捼S�ݖ#�sⶂG^㔅�ƕ����ٸy 3�_4��4eY-��t�\�~)���;wj.{��=��ѩ���yȔ��G��]���)3��+�ȿ3�\�C3Y2��1�E�@�{���9�oÔ�kW�(�,Rm������
�#��#[j!�'��1�.�e�~�;p�?�g���B8_�_%��~S��):��X�S��Z��.�T8�N
����.>����k[ �煍@�ت��l�9��h��J$���J�ˆ���R��;U~xy�v�&�solG��Q/1���s��侼�Lv6��Z����(�q\��
\=F�y�~	ՀJ9��5:��?�P6�:8�Ls,�|��-W�31|��Ù~U���DE�_�+��Q�� �Z�bG��VI��{d��X*�\�ƆV}���'MS��xB����5S�z�=�|���
���t_��G@�5��Ֆ,:�(��uYk	8R#�Վ���b��ԭ�25<�y����ݢ�H/e��/��΍6Kec��,����X1����}l�N���w���z���>��_�ɨE��6l��+p!�Dö���\0�l��}h+��<��'��¼��Q�dR�	¢��rqS_y�����p�xy��b�
%����2�$S����O�i~����K��IN4�+���������I�J��<ٔ{��K ��&�B�>[�	.��Y���^��g�E]J�����1����lP�J�-䳠���	����+6(��8*_&-3b�5��������E3[�)�3���z3u���$~��eU��u���fxb�u,���W�g0&?��G��VI*��@klq��-p�,G����$��d?��Ԁ$!�޿����)?a�cUX{ϖ,t�+�=�w��6�\y�������JAM_�r���Yς�TdȀ�� |)-���B�[����0"��m�A^�5+�+?S�J$��G@�o��pa��1PMg��谌"�j��ԏΫ2�N\��m=>�V�!;�pQ����K-�*�|6y��<���뮖 uh��a�es)��"h�7�1m<�Ñ�-�FߞF`�/8�@�����X��f�����ߕW�x��Ii V)���Y����ξi�w|���V������9���*�L	S���Gy����hBM*�.S������Lp��i�AI�I~N��v�I��%%P<�Q���8v,��v�`6�:
r�Њ$KP	<,��h
61v�/����zL|E�j��H�?�-/��,�*��1.Jf�,R'��W��Jmk��d]|� �bg��'�6��*�̼ڭO;�W�R2,�֧sPvBf���e���Pn-Cr����N��lw�x!��u�KNď�t�yB<�7���O�W�O��%��u����C�	ӄ"����v(��I�)9fL`m�<C�\z����vQuʆ5����.�J�pIPJ��d��≠�ۍj�CC܋S��q������m�lI�
��VJA��xկ�1���E*F���U}��e�[�]��^�q��/��I݀�1���|&_��,I�Q��w
X(��Ÿ�<��Z�Qp6A=>�Dk��b������v�RH��ah
��� ��>��r`��+��Qc��
����2�ۈ�\��r�[�}Z�	H3|4�V��6!Ŀۚ��p����J�{����2�FUID��YƴC�[�>
���ŽV�X"	|��~��V�Xt" n���?z��D���xE�ӻc�ʘ��� �DG$mJ��R�ya=3�v���!:�����O"/�ʼ�m��՛� 7��[���%l�x��w���szD�k�7.p��m,�S�R��Ј�%�[��$�����  ?q��,<��&43��[�4����Ъ�'��/��$T��;��ܳ�µк���H� |��5���]
�H4F:UT��A"[�$���4����6̥�Fy������*-�7��ˏu��m�,��򲨘"0>2���K��T�c� 4�T�e��'S�x�����PC����2[m�y
2BRDp.d��[U6� $�M�/�؅TK.��҄��~��L���C��B�\��ߟ��"����@�c�K�^���0�.��(L��"[7��Au{`J�2U�w�{]or$/,��F���Y2es�A���D�.7���
g�ׄ)��#��"�`�
��p��3�_���R&ە�D���G�`qR���$�I_�����Lߓ�u�0@V��'�,.L]x�����&������"�w =�.����%��"b ��2�֜���?�I��$�����-�������T� 6����("�&r�<}'r�*�-�XFZ�F�V�YJ2���� {��q�5���h&.�Wi" �O��&�V���X+4U2��W�&��N�sO��~���?-Y�%�#���(5Cri��\��t�;$��U{�Jk�b�!�U,��8��9Ģ��B���.��f��$O)w隔Ŝ
��I�"?�YM���'�F�s	�?�d�m�$��Ћ��c�4�ı�����"Ϻ؜��QF�M��u����V$��j�'����i؏y������%��X�����<{H]��l�s�ݑ�c�`�h�"��(;���p�0��T�A���.JbHb����ԫz��%	.��3�'@�F:+��'xQ�v��1�?����ʈ��\_���C*7�|��Zf�j|�8P��m#�o�� �D�?C��O���W��H�հ�D.=�Ӯ�k�l��T�� j��sEI;��O���@��C��XN����8U��AlVؘdW`̟͂#4w��Y@�)d�T���U�kb�\l�{ƖQ{O\��.���ײ���%������S����~���~��?��NՒƁ=.	��N�Ǚ�b��ZR�� X��A�:Ui;� �Χ�ӄ���x��_c�Y�=a���3$0r��%1�y����>�Ra$jR���,p�G6���2v��9%L��A��h�JU�瞄u���:��r5wS�Z~�9b���h7�43�ֹ�i�d�D/3WR��K͖���l��Ѳ��%�#'����U��#h��O�M
)��EI��xɆ�tmw���eb'�<r6�gi������u�͂&�Y��s�4@j�\��u"ء�sA%L;W�d1x�8�����
�a�0�h��/�J0Le�I&B��%N��7��� �;����@L��늕w�2�ݘ��+�&Ƞ���g
PC1��L��b{v�/�~؏Y�ײ�T	$Wr���`�N��.E�Wx%���2����w|@�G*9R�{�����w^I0�ΖϷ1�jP�	���ڔ�򑍲��b���H<�Y�)W��5G^t/Eg)=��Ч�o��Q־�6�ڼ1=��Qm38��}�<�'�5��{4�?g��|�Tr�l�籧�br��D�a���w�hׇ�����B���������v����FY�D��OG�P�y��#\e�J�����~�P�W� �.�pᚂ\��K�I$��'��`���o�"!���#�g�B1议o�t�ͷѢK� ���3T�,n�7����1|��5�H.�eHm�;����2�ȕ#�����۬�ձ�q#YpC�	�M�t_���yOa���!	&0��}����~ZV#���Z*���^{O��Tc�Is��f0��ƌ��K�	b�N[�hKv���M���C�3c�I�=-�X�.t����Ӛ�Q���Q���~��Y_U�d����l�FotY/�[Y��!�r��0�bi�]G5�&��#�Y[k�]��{�[R,�U��v8���=�bDИ���?�跗���:"u@?k4=�X9���I��C6�����7�o`V�<bu3}%-�R��_a���^x'JB��*��ą'_��~Q�d,[�Od�V9=GJ,���X�I�V4x�FV&k�[�$<�Y�F������������������ȍ�I'�.�PI�ƥ��������N��Ѳ�����U=ˣ�+>���l���@~,!]ș���`����{$�����j�n�:�Ø��M�6V%{�xc	��~4L�[�@0CP���L������k�H�bU�ڔ��f����b��T��Ü`" 4�Q�{d�0����h�x��WT��4�ƍ�`�iݣ}���x�J�e�0X��|]��E�R�z�M�T��d�H���<��l��7��t�q��,Ofh�0ij��c�#�' =��
�V��D��[�܎ |#d�O�%�{U��v,�3Fٳo��[m�״�h�2X�9ꯧ����e���N
��͂�=�C�D�CQ����@��Q�F�dBv٥�{70z���le%��pa^�3e>���א86+�;m��1�!,k5+�oﰹε�gb����33N�R�/V����4��B�P��JA�|�I .�ԃ8�����]2}~ԞSm���B�1F�M ����Q��T�������nå'J��*�%ڂ �A=kw��y��՚ Y[I��z��R�?�4l�wK�{��n��S��!2ko�AN!'N��)vU?��B��#ĕ��U9�!L{��t�K~?����]�T�ћ��Z�FT�Ԗ
){gs�a�U���M
�KqI���aŘ�*#��66ԅ*�.��h�b�I�K��={�H�z�ս؎���UG^��~Bl�+�;����:��W@�! 1��(C��\�D��AGZ
��;�CF2�4������&d����wl�Sй4J�l�S	k�S ���yȷ�\����v��9��'K�Y�*&���:'+f���r������$��JLT�K߹k\Y��8v�pω���!�Sc�蚊� ���m�0��A:&�B��$�(�|�-睒�p�tN�9��{"�\:" ,H���踖�<QS�6Ś��>�~�٦|�Y�	��"�X}8����-�xL~�N2���_�1�A"����[A?
����w�����@�c��}��wh����ƺG3=�q�q�T3lX���-�������'м�^t�~��(坲��%��'��L�D����	%O�A*|�
l�r�B��[}��t���ލm4�2����#s7��SFu��S�#�.�I;���$ߚu�ӮӲ����+�D���i�������
�i��U[_)G�-�2�
W\&b6:|-�g�F�ڡ�Xo�Z�nf&{�Y��H}mjy�Z蝡km90�_�C�f$e;�� �y�hV	(y�Lv�Ĳ��BD�!:m�L��,�y��.�����W��� ���5+VL#.�~jC��+fU�����S���K5=Z"��9���@�%�T����Z�g�X7i`����:����fc���O��
�¾�� AX;�ygvz�S�e�3��ZEc���|����u��:i����8A��w����	� ShѡI�� �����7�����z@>��wԕVx%���iV`���B����7v���b�T�]b)	�D`b�*z�� (Uo��l\F���$B��(�xާ*�Z�;K�,`Q��6�a"Q�1逖 �Zi�O��:	�YAu£���Ri���\[Q@KQ��K�,\��%���;�7�I���4���-}\������&=��lb��#6�5_g��w��px���瑊���D�����nn�L2ϴN�L#<a��9lq5�2�P4X���VF2��8�S��Q��E��ο�-.��e��R\M�)H(���mK��� U'�dqO�=N���A��]Ր��|�x��u�w�����Y���X)�@d:�9G�rv�Xv�/���0r�Ƴ�L��IW��88䠾\����/l��i{�<���-[�}��@<����mf��,�.j�����YL�0
��*��?����gZ���'����}��"�,Ɩ�,���'�Z�D�T1Z��3ڛ��+�`d_UTծ����Q4��I[����(r�6n�n�8��n�l��n�cA�����p#�c�~m#�>=�m�}?��f6\Dpp[�P(���0Ռ�0
Z�W��7T��ۏ�d<���8&�!�7:[	���b���f-BC�9`������!����}q��{���s���h�TRd�3"dU�m��I��J��g�LlǖS��.�&u��݂����et|�f)��z���J��Y�W�MmsW,w�X!��m�T~ʟ�����N��c-ouӿG|V�{஋9�W�N�̏��\�0,��K3�M�,��7��=�+�=?w����\�d�J��@w��3�	��S�6M��"��\Ƈ���s�Fv����m#Э#�1�P�3��G'�f�V���%U7��c?�ִf�]HRy�Zj@�(��ˆ������\6t��@�"{��	�p 5u�z疁 +��$��OXy~��ゆ�Л ��M�rf�O�wjH`�F�\��	���	8��H��dq��hc��Cy�K�V��N��X:��e��Ǿ��\��H���[?���Y��=G}�~��7Z�3�Ux�\6��=��lc&�V��4�x���<VF��	y�zXL6+���|FT����y��)� �����:)>X�?9��g�LdP�S!�q�}��fl6xq6���y�oFH�xi���Q�����@ �Q��%�v��@A�q�QrZV�K���XNv	&m}�`��̻��D)�U.M�ɀ۷U�
�0f΂��L��׃.g{"PC�/��='���q�a8��&�eiӥE��]��M���kQ}�E���tī���1-���R�Dpv���M�Df�M��؆`ҭE
І)�����E��j=�P�?�	=�-���G6f)↤���]�&6����䷾����$�<���c�4�(�c�>?� :���y	"O��;�v��yYYL/`u��b���.nqp����Wj�
�HB�E�Y��ѿ���!�I��*�Ꙟy7jBs�h�;,��ԅH�!pf���E�|�JP�W����q2+�~�ھu1�$U�Zi��k���M��^F��h'�t1�G���떾���1����$.�<����.x%jؒ�C����t��!LĿG���Ñ������n�����UES֖�Cq-�n�Bʛ-P1̠��yϘ�+�֎�]u��fD1ZIT��Q�z��1�/2m����_�Sb�7ˡ�꺤A���J���)h��K딷{+M�/��e�H��<�^����N�����U��tdŶ�f�%HP$��p�R�5Z�<����8>KoW|+�A���L-;y-�6��K�i����"e�J�.�J*�JMË\~-��.2�ߍ��n�F[��Z����o��Ճ��v$���4٫ R˭^�l�k�1u�����
 �ޘ"NMh����Wp��B��r�h�5&I;�"򐇓!j�3yfv�W�DX�4s�61C�\?#'V4څ�qM��-nÎ���թ��2��r��B'�~����Ē�������B�i��&�a�ǯ�a�	�H�߰�����eHe�ǧ���Tb�pf[���)[KO�,a/jmw�Gܤ�3i��UрS�%H��S[�����-��P�l�Sg=����It)s�{c�[��� �:�x��^�Si"u�az71� �&��>sV�2��}�륈4U��I��
�����P�c���������m��hl�����1���imp��$��E�a���Q!���Ƹl��n5��h���:����d��C�xj�+���!`�σ(�`��y�V�t�B$�G��5����;��p��8;���s��4�23�������Fn8?
�2��c��8���V�*fh����^?}�"�B����͛C��s�����]Os^Io%n]N���O+m���-8]3긒���j$���g�s�0z�j�Y��+�o����e��}���鰶�	
�����_q���T>�&.Ѣ�H�D����9����4H��0�0$��%g ׶�K��`C,��c�]��U��X&)��S<��R�X6�I�L�㙸�ː�l].l��0�W�kD��I[w�������X�єu�)�2�v�����)Ѥ��R� �D
���9��uA}R~�ݑ�AR��Sw��&��aH����e��&�0?y�7y0D��0��n9]l��#)͹�����tG������P�D�)�n��>�{�Pu�ᙼ�^l|Th�q�D�$������
x	��W_���e���Θ�]]���r9W�±Y��mif9|�5��`�i�&�8a�L��u��&�T,���$��M��ϛ;����-y��:C�'��?nT�[�5�6�3���R,nyBޛF�_��љ[�O\x���EH��tS�A��ct��Y�� ���9U��\�e�_^µ�¥�,��v��C�~�P�o��-�I��`ހ�Ig�ت I�۽�T�Hg�"S{�����3?�G�	}Im�G�{�9���i���bjc<s6mǤ��`Ѭr�{!z�[�Hv1h@~6�m��D�跴2��<r@��,Geu0��-`m�~
d+���ⷭo���.����s�3���a�Qn����o{��(:c"9`%�ޙ���7$����
�
�:|�`(QF �������e"/���a�מ9@�w�ܦ�h4����ڰ��O�	I2���(�6���#uQ8�d��J�Ki���nA��@���su�"TL(;R�ݎ�t�I�G����1a�R�ɮ|#N]!��6��f��N-��Gv��U5*�8���#�vo��EPA�a�q�`��2Aб�e\�sZ�_jԘsră�� �].0l���ɏ��	�e����a3�K�˾��2f-���l�˧�ɻ#�7.�G��+�D�;Ը$7�U;<�v��(�~�P ��2��~"M�*F�İ�W�J�٢��ןu�I�Æ:@[�~n�ʁs�[L~��ٞ����p6�x������E5\ܐ�rO�<��غ�("Z�hqC��ݙغ�@g⋵��4��]l(�(%�aR�r�6>���{�.b�8�8e���y�M|��~�	��$�`x���C�.x��o��ж8�I��ek�j*��������)�-�������!��v��y>Cn�b=�f�2�_���Gi�K����M�^�>��f"����"=S�tNk�m��)7��c�ˡg���|?�!�L�+�Wlq|Gܳ��R
��n�t�ƌ/����^6в��nE�>Y����xR@ڮUԩ��x5�̳4q�c.,v��گ���+��+�?�Oc�� ��}�Fښ�u �MmT!����_M�;���?���_�tFi^�m��w�U��6CӪ��p�	>ڀ;�d`�����7ȯ�5�V��&û�\��$�}�\� *F�t�x��;��Ew�P��W�^� �~W���Qq#{]�7�2=-�9��(3�-��
R%� 
���qV<��q�c�{8�/^�%^D_���+c�
>�}�Y*�[�����kh�J��V���Q��*�xh�P�!�$��;�����hW�劇�+��Rhhc����R��ÐKɿd����G:�^��,d����}yI�آ\�Wx���2�gvF%��?�-�ţ4�#��ht�ҰH����>��`G�+V�`�a�O$��ep�{,wd ��K/?t�dG����ձs��H`���F�*Ț��\�?)U�������f�EÿZI��٭��é���-�X {dx���ظi����������f�f(H�Ep+M��P(�9%lD�|*4T���ڳ�x�ֱ!�V�u�ܢ6���D��e�͞�F�B�Bj�'�&:�� �a��h��4��Ⓛ����L.E�;����97O>-��rq=+�������1��1��5Я�q�7�����38���Pr��[�w�هI�?���I��)irY�:�P,��KZ&@��z����7Edu��r=�T{u��l�͑���_�5�}!�c�r��cٿ�>���L����y٬C���������#"�kԑ�[:e�*��[e��wJ����J(��A�'��z>1Q��'="ʴ�@Q, '߾�?��("أs��7�$��B�*�-���%��э��9R�\'�>�9�T[��o�c��C��S_R�\E���UH�%#���;��&uܭ�X&m�+j�<�8�,��l�'���F*'�W��s��̩MK�OU+���Ezj��N%dk��
y�������S����È	���Y���~��E{<y��>�R�D�%z��˹*췾�� Y����:/(s�+䵛��r�)ۄ��qW���Om� ���Ri���1����P#�ur2�U�_�A�y������}M5ѻ�:�߹�+�_� �΄�T1��o?�K�����z��A����[y�r����ç
|���!�]�����4�8���R۬�FKK��8��9����=gS�";�;�"r�D�{eJ�P��i���B�Az�$����d�tӶ�8�����j��cR���ߟ��os��C����
g�
�>2�I��A���p��l�g����V���#�3Ζ'm��]ZȰAS��
M�F��$�O��IƢ.s��k�����<�eaT��Q�C�!e@��ĸ�h<&�8��R�,ʔ��Fr���@o_�Ed�~��	Ǻ���yɷ6Ȗf�3�1�l���LiI1)2�4]W�-9���L�L7�^GGN�H��Po��&C#~Z�2�O9�%�yӱ��X�X����N�x!��G�@fI�C�̩�Z�am�� �K��ʂ)
o�����3Id���b����r$��6�w���e�(:��0hM��a�9��q�?�d2^aD�l�Ps�Z�Z�\����R�a�z��"��
��K{�( /p�?�]�������G\O����|:�6VD?��T�k��z���7���z���,ph#x4r3�t
Z�9j��y.C<���S��s���U�U�_6�h�9��a�M�j�0|w��(n[9���Q�Pr���hD������:z��K��o�8����(�jn��ڵ�����⓰�r���I�yyi �>�F JF��V�R���!���%"�0ϡm��.��3;�#q�d#��W�i������V9��v���3��)#�p�Z�j�y�������yN#���w�KH����.�vl�*X�&����Z̊Z��pWC|@���5�4�w�%���J��X�s�<IIR�ߘ��N9�
�����)��s��m�]6��w���@�v(���M���|rN��Uz'����#aTMՑy,�|�I|Y1�8��(���� V�Ha�ܬ�?�F[�[2 U�����C��<g�v����b�#�B�.��G��a,^q	���A�G �j���v��������b���3�W�3V��,���"�~��+�P���黰.�E���:v�|���y�� �C��u���@��sv3z�^���|��M��,���g �޸_8��5�:[1�#e�>��*��K��cO�zs�P��@h�<���dS�^�M�-s�T>fؑi�%"� ���j�	�G���3/mpF�^�^޵n�g�M�`��� ��8�_O�5���i�A�E���vwP���I�|z��4�ޭ�Bz��B2�P,'HG��:�5�z�p���Q��k)�bZjY�W�����:hR`E��IP"���;Z7��f�te������w�\�<\����_�+F�+��S�Y^��a��s$}4�#�A�����7���>�iMa�b�o�+0rCG_h>���yh�_Q��5Ǔ�3�Z��J�c��7q��r�B<ȃY�l��.s�È3=���n��;�
9������$�()D6'�p��:�W����a�Rp=:5`x�=@�̷/�Dq_t��V�0���zh�k��i���v!u�b�^��3���Z��k��PU�L\���:
�t�=�)��p�w�f3��'5��9��&5���e;�uKme���2����� ���~��@؝rי��#�[w30]
a�PK5��[��_��S��;P�"cf�e|�j@�Up��4�ZdWL�[$��{O�"�������F�����������~�UD�%}SI�����jK��8Z	����֪1o���_8f�ρ����JJ����; �/����;����Ə�,|@��L��A�?�N�� ,~}?^��5vb��*I��㭆����|�f PI��S%�|Y��;xz��������w�uen�c�X�9�}���~�oc��-�Ԅa;d�e�4�jY������ț�m�g�kKı���{�zlGn)m�_rq/A�R���ht�\8�&S+�d�Va+0s/;�#@���C�]�x��J7���ܪtB�Qv L��oi��΂+	�Wb��8Y'���Sz/(���Š.��	f �z��|,)Q��^P�:���ipa�ￎ�}��6v�ǖӜ�ncV��R&�-�5t���(߂K�A�M/�P��*֒!m����;X�C���Kh��,Z��_�+BfR�:��� 5���I���,�0E' Kq̈́��4�/�{���97�g0(kG�e�}���gf°*��`���B2�m���Y|>��݊��W�~�m�M<?�'XV����+�L:�V�|!ܘKz�*ld���.}�������:���g&��q�-�P���V��Đ�m=k�)����'�s��Ԍ�zkI4�{F����0��FS�R�������4��Q���M�"�0�QQ� ���������8��u�=�t��\��.ͫ��NJ��W�5�q?w&7yD��%�
m;��ot��ue<�v���s��A�9�.�)�C�����ŘFZ�D��\y�������2�yԘ:2CS��>��=��c&y� ���	G�3�Kw.�̝;9&��L"
 �S9���~~g��{����e�|�-�"[۬҇�b�Գ���zWn.1d�J)C�j��0BD�fi�{���P��ܰy���H��	
���ڮ��\�':�[Q��5�s4�$k��K���]��(� l[�SQ�O]��E�Ե'j�	���Ƣ\z�/M���@�2�E
`�����k��o�}�(��M���?˼o�����.a��k�Ȯ�%�_��&A^ 6���S����2o=Z� ��-S����۝1x7=Y� FH������E�`��a�˄�a%�*��Hi�m\�>�o����&ۺ"ڏ��A�������q�4e��3���Z1=����_�����:7�9�������0P�&�48#��	�ޢ$��|iKK��t'D���\�r��r��g�&6�+�#���S�!�ተ������'���X�j�td�rW�������Ϙ&�`ԗ�&!
:�q`C#!M$MX�]��:�b9R"�/Z6�9�
�*�� n�?,k�/�g� GCL�\S{�"K떰\�i�s�9H�<9�j�f2�뛁�B\�il�3A���󪝂���a3i[�K2&&�#N?��p�z�6X�e��&Y�3{Y�慻
yµ�Ԓ�	�`a��`ડ�Q�u���^V ��SF�����~"W{���0g�Y�u��?�6��C�+nC`d^"�9����)�"ɸ���o-̝��,�k��M�Z@RX�"�*����-�E' uT�QX��P�{2-�[���΋Ԑۯ���7SFq^8��]<1��"#���1��L�΀���Zw/u/R��r�v��>OL�bWR~�x� ����Ww��n�S�td<��#Rr/A�+�&���	8�H�B�`���_�Ƴ�f�s3$�ǂY��M�. `J-!Z�.鄑{��o#��@�������8���S8�~����b�����*�;���?���M6+�5q��G�-]QV���%On<��~��*�o��9��&�\�d�e{0��<]���ȶ"Y|u"�m2I�lh��Z��2B�mg��ɳ+�_�OnB�D��Q�fɱ���r��k�U h7��c��bnO�p�,vV/*%v/k��Di��Ү>6�F�Q�*:\XcNp\A���w����uϧ�	l,�0u�@`۵�*1��X��Bj�����ܬ1F](!k�A�Rb��4�鄁V���3p�Z
6�a8`���$��T���w/�U��/]��=��/<�Ic-yf�P��_?`p+M @�M�e�Mw�ޤa�	T����u�#5[3p�A�ܑGM]�"v�X�Wka�W�X#F��~�������.L%�Ԅ�x78��&�!���e���.�a	1��hI\���x���d�q~�p��iS*X��,@��X�C��$�C!jj?�����- �DhW���=>���bx����_#4 _)	߀+ͅ�~���J�psf�C=�D�ٖ
�ϬO�rd�!l�O��_U%^���d�����7�Aw������6�=. �CF'�����#pQG���"�F���J�yc��^b
x�;���лW[��Çފ�sʦ�m�!"�E��>֊Hy�HJ$O�='V�k?�
��cn�n�DTE��~p��t=�9�շc���u���WJ��c҈+�[��_����9y�w�/��\{ٺ`�m/�`P\�'h2� �Qh��Hh'_w�ȽL�S��Р����_"�l�4vD�A�*r`��S������lG��'�iz�����'��Gk��+�E�
�g�<��FI��� �dL<M\zTV�v�����e`��>�k�tI�)e}|RN��4��d:_u.�i��D�j�G�[���y5�q�a�T�;MelDad1�����p�6�f`u��3�vE�m����*�)3�U0�ԿRO�譆�!O�be�m��]�	)Ӿ'�/�3(Ɥs�4��k��5�b��8��)!$�����K|�>
uK�Y�g�ݾ���b���f�dON�������k���8R����O��T�7pUp$~���{��x��bR��c�Ӱ��<vAa��/�)?��p��B�Ui~U1�"��|��%�M�J^� ��/���x|z���{��$���2!�20��hL�����S������0X[�!D*���+��,�0,�t)Dⵦ��Φ�=�Єs%�h������1`Q؏~آ��#I��5Z8���9՝4T%��',�8G<u�l?�{9�ʐ����Zz�a�/N�����/��2NFTE���NiA56���Q@�pHk��]�+����[Az܉\���(��� ��d�`uk�>9Y�bMԎ��J���D����.-����猽�坠�ѻED����ğ�ilk�k��}�;5�L�Q~cI'���=�w�jt���r�������Yi'�5M`�,R���L�8Io=��`�O+57��4}�-������}��n�.�-��y)�3��Ӓ����k�r2w�鍅#v�?���)9�O�����)����HI��K~o�K��Ǝ1��֔��vk�!��N&��،Fǵ�n���B�^��n�7+���Ц0�u�:��!6�>�Aij�X"��pr�Ԙ'ғ\�p�d����!��8D��Z��n�0c�?����Rfq�L����W�ao7o�c��:8� Uj|�𚾷��t&YD�߅]-��V/x*���Q��4�w���{ ,����|��f���?�V��AE���v��S�E�l��/�?��Ҕ^���Λ~��(�׳�da�*�_��˰b R�`���q�P�x�gӛR�U$	BF;A7�0�'.��@\lza�վ��ĝ��1�hYT�րM�AI1��0h}����5Arl��v�'1�|�Nr����X�#�����zs3��2��\vF��x�8a��)���/<O�+�@Zr�D���񱒳��H(f��5^�ЦE���e�<�b=TV�� ]�ߗi�����G{��TEB��|�[�ñ{�r�ⷿ�ےT��˴̼_�<�'�����P<u�KB���,s�S�%���\Y.��B^�^�����N|�}��Y�G��ٻ�х�f���v�b҂4z1�!R�Iբ�ꜛ.8��P��J1�b�������lS�E�ˎT%��9J�*]�j7'%�UP�?+�S��l+�*�!�i"J�S��T���WL+�PE��L=��u�`�����|���
υ�b)-%N900Qi�Q���a�fÛ��#E���ݘ��c	�V�d��P���"�D�]Ԟ	1\�
�/��&asLW\�M+��Qg'2�����u�
�?qp���F9��Z���7�Iɑ���|\���*�H �+s������taw���G/A���9�ŭ���p��q���B11H��zy�"�r<JP���&FI~8�@NOm�y�t�]�Zqz���0��sOtc�����	sZ�K섥��pgb���ʊ�����dv�fL*�cl��\��D��ɢ�,���R�C�E�F�n�Ʈ�%�C���V2e�s�{j�}�Q�V �ȒF����	�qs9]�J���0bQ�{zq:��U�hϘ14c^V���%���(�[���ͫ{�i��ڂRW~��.���������V$�D���� TwA"�4��^$Ys�%c%�|��h�h�Bɮ�����sh�оѡn^���4D��֙�ܠ���� ��\l����|_��6���[�1��p��5H���~^��K&�T�>�~M���-]��e���!ٛG)?�N!#��h�d�inH�B�Ԟ�?��@UC��^��5����f�	�u��J.>:�-���e��1v��o�j&�W��M��I=� ����"��xN�]��Wy/L-n۝a����C!�XƐ�n(�s~&����_�M �Ԁ��J���MVS���t��yZk��*<���'e.G�1z�9�Ѷ���A�o��\}H�g����� i���]b�IA:���>�G�\m_e�t�5�w�q(Q�WnW-�l�8R2ͥ};Z��,��P��pEJѳ�����-�)�)�C���Z���`��S�ѮH 4l��uP��;k�CI�KbJ��"��/�6�	�V�W��f�Y)�w~V�']��fj��\"=j�iU�vr�C��23��g"��<n�OL}VNh��!p�]�T�D��#�L&|+?�^^�#���Ǔąr�*�����li.&�vt��+\�S��Ǹ��o�K<Њ��Տ��.mp� �]��ĺ�7Ɯ���\U+p�W>:�q��}�� �
�Z��4��5��Х�q��` ��t��
ve��z��� e6�$�uL���[�@!�&+�v�SE�y�n��u�7t���|�gn��?d�uP^;1H&.�|�Y��|֣ ��_%J��$كKM���syKN��h(�n�x���C���sC�f������T)fa�$!N?<��ј���H���5�m,�ɭ��{/|fm�a�Q�vGF�)��sv�|�{�>�u�����^�#/�5U'
���_�o� ?"J�{m�^'�k�(4 �n����mX	�|5���K�������op�,܅t�K��]g��j�4��8| ����Y٢��D%V�|���<<��w�JM��׷��ƴ��߼פ#$n�+f'	k~K���Mw�=�"Tm�K@�fb �R-�1K"��_�`K�%�)I�f����1b�1�r<
X���z� �����n)U��ò����WE�Cya���eS�-]����U$B���}NLٙ2C���-2~轋�f*�?�^zQ��r��[.���[^:c/ ��J���=�)a�D*�s4d������}t��pR ��Y-Z��3��:��@1P|���	�er���hQt�Y�;X"x�aC<�7���ߕr�qмѺ;p.����gX�Z�o�q�y�}.���&�0��0�³�c�§�g:,0�G�+������^SC�ʭJt���!����+�3)�x��|��N���Ҕ!�.U�������.�t�� ��;���nM'j"�����A�5��H|�t/��E��*����Qkr��vy�+�,zo���sZ���Iʇ���%|v��%��"<��O&�JKն�(�wɗ�uX"�$g�~���C�/T�o�
�~�(l- �Eioz��P���O}��UӺ7ǙdY�Iĸ���%��Z��:SX#�^�����E�f�x�I�d�d�k��K��K§�4݃��$��b�u�л7����_��	�hM�>r&f��/���۴7S���t&)ퟥ�L�q�x��aF��N�MG�g�� �|��f��G�P:���9��u�{�-3����2��U	��z4;��jo�1�B̽���6ڗlbL�-G�����-=о�g��ͬ�-a��������|zLJ�0'��Q��QM?��^��(O	� ��˦KoL:HJ��[��K�d[���J�H��k_�I�I�����͜TA.���9X~11.��C��:���j%�M5Wd8��9M�����;�̝���<�t����k��a��]�ɂ��� �bK�̺�{?FsW�����	F[UI ����`j6wE�#��.����=q_#]��K��^)l�A*=��g���5�͝��A�0\�]+��?ўd
y�h�S�8�@ ^�����"i� �+H������
ҝ����	 �)^]��]n�7	���7�������w��1�y��:x�lǜSfó����a��=�E�AyE�آ���Ď�p�������͟.�Uv���^��|\��坴�k��)cC��"|e���ʑT6}�̓����%^�D���9f(��%VG-�gd��AXYYȓ�r��Mv�_��n�$�j�x��X6$�]*��<7!6T���\,���3��4S����S��\ Sha�`���.7��L��F֩��%;��$�9��
����E�F����l�)�pTֻ3u� �5�V5��]ҢJGr�aY'A�
VZ��g��Z�A�9���+����e>�,	�h=E���<���]~D�f�O�M�t���e�u�"�L�6Il��B�]��a��Mz/�B Tc��iw,��r�ɛ���U����JPBw�(�;�?f�t)��=h<�Y�XS�+���`�w���55J�q�yQ����d��悗m��$�J��s�TѨ/\l��ۧ+�J�� �R��{�8�`�0��gh��"l�=K�j�,�0�V_�YI��'�X*E�ȯ����:+�]�x!+�*���ǂ���i+���]3��R�L��C;���Un���S�81�A�>1�+��$~�	+��Տ����j����(�������#�|ؘ[e�-S��U�1d5VE��G��69�L�����4���}x���Jt=CS2��ii��{#sQ�n���J�h�hw��_[���v��^XsW]z>�{�0���"�/�~������c0H�L�}��R�N�Z[���2� 
�Z�'|StV��Vb�����G��0�ےn�ިᔙ���4�I�'������4�e-�5��(���1�̮s�ZX^��ݐ�嚄aq9���q�0#0�t��벬�;�MN��A�Uu�9͢O�ӕ���@׆Upxvpzo��7�61���`����;����^��n�pi�I-LEYh�yb�󠠚��?s�c��x�@�^���Q(z������� �g93��+����<����A!v|(7S�n�����o��xmP�,�X\�C�fF��a���~��%R)4�{YE��V����"{�G�;���:������v(:8R���>�F��Z�
�q%w83���Y��ꈩY4F����y�Ԉs�B�%��WlX���V�����O�k��{�v,!��j���qh�Ʒ��x'
]�-��3�ʝѐ*�DI[�e���þqS(N=���>��5<vU ���DyL���������f���QU�)�x�~�7G� �c�^�r�;~u"+g_2�Y�[9hJ���Mq�2u0��k�a�,c�h�Eni��� uC9��'����4�%��5�?�AN�@Vj�ì۴�Փ��n�]�AB���J%|��wS6EVX���>�e�D�`�X�VY��/k�aq)r��=7�F��.���â4U������ �0� C��TfLQ9`F�������^'�X�6�A3�����%�v�Yǅ�<W�[�Vv���.;g���^�@ď�Λ�y�D��m���o�:{mG��ݏa񯓝�������%�������Fc�����c'�R�򗩌�:�z�� ���X
;�"-�T;9�B�.���ɶa��#Kjh(yn0ݏ��1y��5B���5�a(�����]&��.�H�#�y�[���;�~��/�X�n̢X%���`�y� 
Q�{�և��ϥC� ��c�x(�|(�$.�B+N[_XDh�� �ء��2#�`�|������)�S��xk���H5��x���nh�}.ʔͭN�~�5���!F�!�-��5�6�V��0�B�3
Pjj$�6~iӋ��z߻��C���3[������m )�;5qa&��2��|!���b%��ޤ���l<��3���hQJ�2�o��?�&zw�&�Z�ji���u�n��9�_d��OO�R�ޣ{A�@���yg(if���$��]���=ay��$y	�>��j1:i�ci�k�k%|	6����J�r�)�~�����!����W��5�SV�i���{3�1��}]<�$u"�t([i��֬YDk��
}�Ȃ�#IG��m��v���`|�������g��S5]�歄E�ZQi�;�K�Ű�,��+f��1�B]v�+,t�,� �'�k���$��#˄��&]:2���7�.�.)O���7G�	�e�c�O�]zm�ζ�u�B`�rA��"7�	����1���Q�ڗ`�����%���� ��u.��x{�K��V��=����ގ����}�~H?j`�t�8�Ʈ.}
��m�NZ���ӒXg����w�4�c7$��\fXg��'Z�+�`p&@�2��%���c
֨��Lu):K�?d9`Cz�G-��}��?�/
��ud��Wu>ۇG�B!QDD[�/*&��Ǯ��#�Zf�)���'>�M� ��ַ�j�ư���o��������p:~=KF,r���Ȓg3��/�%�,�r|-��k����~�\�$�{��w�����j��X��K�E�"�JV��Ȗ�ؿ���%������o���k���I9�-2��u�{o�x'�֎�n6������Ͽ)̃��ݰu��߆��g��I����<
�0�өŮ������q8%
g���$���w]!%�/��Y'�F�!$� �2;�9�h�nAZ�]��C������e��ߚ{d�I�-�u�i9�-e�)�J�SO�\��vâԉp�p��uI�3oe�M�D����v��<��h G��ێǕ�ue[����+������Oȟ�E������'K�C��BD�5���?� %�䃛#���c��mNG��\df/Z����XbI<�;e�#�A��Ot�P-[�kS�`�w����~��n� �78Q��ǪB�Rn�^�b�ml�
�P)����?Z`t����P���A�l] �Bއh)և��[a�.�Vakl&��Ɩm�4�� ����e�n�Xr��
{Z�A��*̺?�W�S���NGc�'q��k���꧊Ca+�-`��e�ҞSRS@��*`NGd��G�M��9v��oD��,�2A���ǊݸՊr�Σ��a��<���1���(�	|{�-��@�AW�ʸg�gx���}FƏ\Q��*!ǐk�˕����'���s:�z:eP�Gx.\_�hp�o��
���}�Ʋ��0���24�������ѳr:����sHTQz擘_̊�R���B�;�����(B^������oR���/i����
j��~ubb�#k��ʈ�Mo�q3����k�tc2����,c������#0):'n��CoX;��b�j"�C�%RH������F��0�/jW���C����B�*Rߜ�ny+bi�-��]Bn���F�O���1�(7K���Z��;�g��Z�(Gq��b�JT�b��]5I�s��A�җ@��(�(�uM�)�4Uy�^�%ӂ^k��{2�u�
�(!������5RmR�e1ZJ"K�@Ҭx�eͬ������6 ��w�Z�D�H#MW����\z��2��~��Y:D�V[UT�^]ؙ(w�3�s��gVObk��=c�2�P�;w��2�o%���E��SL��C�swj!H���þ��Gf���Q:��y	4�%#D�5P"�x+�
�Uy�O��޴m딑����e$�{���7�6KQ��״T󲣥��'�$ �(9���*C���柬��MN��f���fu��t��M;x��*h˜�}@�q��u	�z}�j�1y�,W��ε�8c���#h���j���z<�46>8�;Βw�B��E���������@��D0������z���{��O� ��c��W:���.�w���`��S*�����������o���2�ŤD=�!;��8����P�W�9-���S:�����I�m&��EX�pi�tu�̌���z��R�����x��+jo�S�P�������{A���7���;Twțŝ�'�a�2i���rA\���0���, (\:��d߽w�v�ҽ
@�~��A��F��UT��Y�s/@q�ԥV��vCϏ�a�A�����0��-��0ܑ�H��{j��3�Vݣ."��u�M��F�k1:�8��n.ҏ��@L�����'��;������=B�i�zzG=�MJ2
i�<��r�CR��pSĸ�-'j&b&N�E�Ϻ��Aq2��o���#��[��m	�zJ��l��>Ge����8g��t�"q�((���\C�idk{jGn��(��=�G YS1�h�~g��We#��72��k���1=L�C�xW3�0��B�kTq��4A'���~TvkX��|�B>��>�*#��9���>
�Dc��7Kyʞ%.J����v�i�A��6U$m�7�Ơ����ryĎxS��[F����e����Au�h��Gǈ9�� -�\�)Q� |PN�*\���O�����}">��؉�;�-I��
����Vk@��̩�$@��Dĵ2�C�@)����M��2���5ҽ,�LB�'0��X�LB`P�eG��wאL��(��|�r�N��d���|���v�mW6�R՗�e�52��!��N�����<	��!t;�C/M��x�� ���_�R=t�7~�=|� [;�UI��l��"b?��o쐐͛�-Ԉ�� .��5%�`�Ax	|�
u*����u]_�#���B�?ʡ*���3*�o��(~�ק%�!��hˮ�X���ѝot]<m�5{1w���z���C�s��a�j�� aEA�5S����٥R�H#g��V������{��G�H���*��
s�x,���Zdȷ���|��	$ֲ�)�x{KŴ��Z�2���Ւ����S"� ٓ8p�o��s�=ȟ���j������*�|��Q���S���b��q&�L�W׏�����{!Rɻ��$�%\q�2<iΣy��85	���f@&�R?� �ՀA�I:o�Nu�qI�����7B�a��P�G��@���QE��7V�X�Q���*q_Տa�,�Њ]r��Z����j�Z"-'z���ȏ����!c}a��Fj>��~V��=�ѬE�$���9D������k����W�ex����|-�o�lg������擦����������fQCX���0�0������8\b�!�=p:,fF�v�x������̸��5�c����q§v^T��*�c��-h��O���Ҋnُ�'.�f��t?���C�d�L��?g�?�ԯ@5g����0p�l#漽+N��w���c��ļ��ПgK�ky�o��j'%p���o|�P���CKWZf�=-.-��F5B�oN��o����}*�lW��ۮIWE��PA�=F��BjuK&�!�mJ`��efƑ�0/�~$�K�@��ͺ����D�p�T��WL�x<&�c:��t�]���.����,�+_(�����������?�@���}(2	�Ϳ�P���X�&���&��	�+pp����ɛfno�y��'��v��_������F��a[����nn�Q�^�Ő���i�l���D�5ݜt�PD�vGL�C7�.Q\sU�|eC'Z�8$���>���,*��wdjrX&yV��X�T��X?�qn�&M�S j[?�q=[���-q�������B/��@="�z �����}�"?F��qq��p'	���$�v@��"ëyr�1����:�[1�+�Ș�u=�,��ۚӚ�~V!�����Q�)w�0Y�H��i��������~���ycc�1vd�m�|b4_���ỏ~pp{�RU�xl6Z&�H��"h������6,Q8�u��)W���XW�*��Fs�S˻�%�H�_�}6C>q�\��6�{9��tYXY5/N*1ЧpPi:���\���S�z�&Mx�O�Ɯ"q/������^��k�y� ���9E���x�������Q��"���a��]�傒�OzT2���k"����l�(�o��b�嫗ZVKv=?۲����`M2�N�00Դ���OSI7�W@ �p��C�;N dY��9^oi�s}UY4U)&�u�U�߁��y��Ne[�3���Q��:%���K��nK"U��W�:!���H�5�8'@�B�?��3Gs}��3�sH9����w`�U�/;���+�>�ʲ��;n�Ȕ�Jq��I����Nk����
���
Ұ�����D&*�	k��v܏r"h{/��E��zM��>�ז�Y�ǩ�G2;&+��6�1=�ƨӬ���O�o�&
#~������:��e��$�>�c'"L��f=��#���@ڹ[}���즟��'N��ד��������%�n�1N����Jrw�f���A�;v�z�ѧ������-#��%����K��QCi��U�-�uV��G0���Q�O�9£%�pk�aD1{Vn��rs�j��f8���N�����C�����ұ;O	X��(k;]:%�+4�Q��JoF�[�{�\��\�j��!��3��X!4t�IʹDjf~������N���5x��;/�b<���kv�w�BNE��SQ4�W 򑝫
g�  bu�1�W76,�����Tg�}��Oq���/�����w�x ���}LyS9u��t�/0&��n8�e�!H/�u��Q���k��0+�4=�̷�\�� ��bf����q�������MViw��>(Tjy�$�LO窥Q!c�y��S��ˈ@�sXi�lj�U,�V��}��r���W����� ��m��&�z�-�&�@?O�g9����U�6��	��~�ʯ�<u#�86���@�+�`���hVp�41� ���u�y���4�0Vw�U\h��;��Ŝ9��x�~���SO��CZ�*�ɌQ?�3�<����rWb�7��}	丁 hI�,��vm]=n�;�m���f��Ֆ���h1|3Lf�k�hX��y>�7�{俜YB�"�6�6} �K	�}�)�Of}�S�P��������c��r�P\㵽٧���j]
}^G2�,���X�9��ڴ��[�������6^�=J���K[M�������QĠ<�e����i��lyV��T����s��k���R./sH9V�H��_�_ёf��mv��=����c���_���xdH�r痿~e�݀���3��<lp�*��#N"�-E�����8���D��U�c:B�ߘOl���bW�w~���4]&v�=~})�4��F�ڤ����$�9#��s�ti��Ay��z�V�pb�
�����(���Ƅnu���m�?t�#����㕰���(�t}��F�\��6h�1��p'd@�q+��7bq�?=�"���`p[�������:Y�#ZJ,֟�h|"z�I��m�_g�w��~C<H��V*nVk@]�t��\��cU����E}:�&5�29u���Jm���M5�;�Y��F��X!]��7�.~�O�H퇤��S��J�.��=����EG�Ts˸�Q��/kVW�j���Ϝ��ƪ<�a�Q��r3��F�[�C6:z%+���\rx���3����L��S��dC�X	��|#�4���)99�#��O!�u��f�CQ~`T��aJ+���"�s;��mi˯��ʇ���Gh�"�6�n�1h��d�Z�
	 ��\mhil�6�����n�Tޅ2�:��_��C~7v��y>�䐟�tg�S���g���'Nu�o��N[m�_�Mt�>s�A��"��VQ�6�C����$� ڢf��ƙ���::s���Yj��;<Yо���ԫ-M���~���K�a��,��l����[����Æ��ُ��q*�����pr���t�N���Oze��1H������1��)y^��x9�7�,ʒ�X�˙�@��޽�.o�2=}Iv����r	$&Ki{�$�\��p��_R�|��![[���?�]z�F�y�7��[��z�H�����+,�5D��o/���y<���O��=Sj�]{�nX�}���qQ~.�L)�J+|Y��%�3%�_�Pv�F����еt�2Oī����N�2m�iݙ������n�	pVLo�����;y�ĝ'�ֹT��_� #��*��J�w�PwTO�s��w����࿼�H^#�KW��m0<�A�[f> �Z��w�g��|z�sh����]�}��P�vda�e��[M�P`q~�c$*��b&�A|?\-�z��bWwųe��O��׍���Pd%c�B���S��skx)��0C�NG�|**�.�8v������g��w����g�������� �g@�8|{����ՙ
��]U�a
��#J
g,�V?K����p���ݵ*o{I_O36�Վv
�@�~k� �TZR��s��p�m��&"]���Y�7PB��&��6�#aS�$8����)( ]mmHv�$��� 醃��EF�%I?��AH�S����湐�C�Xjǿ1�e� h����i5�����*s�K�}���$��F8
?b����4O/m�s�O�2Lb��QQ��X'������~���Ѿv�P����h���Cl.1I���Ņ��k7�4ԯ'�f�z�1�W�(�l���g�3�*����ډe5��miYjd9��qB���5,�-�qVZ��R�5P�s����WeY؉:Ro�ԡ7.X��b��h���W{CQE��҂2����eQ'���H9��J(�X�_����N�``�I�#k���(�Ψ��>�K;��9�kBc^����� ���5��\;ׯbլ��%#��=���!��j�� -z/by>li�ǐ���`ے����r�l��~�l�g%������;,4f	�Y����|��$����� m�w�d�@�@�7���0ו��J�R���>O�
��Y[�}+�}�?���UZ��HހO_��]�_˸w�N7a���Ns��A�d�rYi	��\Z�~'�	��B-<�Ma彴H*''�L����X&�s��T�5��:�c"�%�@���e���Bb���n�H�"����)찪M3�9�m����є�5�?Lo���2��81��mW��%�{OWQ�;�r����QA�ƫ:���7B�6�W�T�)���B�hY%z'��J�}��V��+�fyk�@1S���$�	z�!�Jbm�����[�Cv���Rd�F��J �x�l����4���<�x�J����^j<p��<g<Ԫ0� �Gկ�v_�`��+���KkH����e&뼶'Wb=(�H��FđE9��3�����=�����/��j�G���%��5��3����Ԑ�.���UDi������fÓ�w��]��<��=�����;����O*|SPg��DJ ��c�w���l���y@

��y�����i�xt*`�G��3ds���<����NZ҉�G'��4�#�q�]͉�������¸1	����߯�}06W�ٟ�fIv�B�^�=` �!��T �S>��|9_n�������
��  ��
M�<�eS%n����8;��f�����ݘ��(�����*��qdY�`�,k�ڽ��0�>�v�5��9�v���G����ER�dcC.�?�s��A�-�r�s+5��ւ�-P�U�:(��g����Q���D����}�R�Z�q�,�9#�,VN�=ܹ�tBׯ˿9�G55}�(�v���ߑ���(F��#��n\��A~�lupx���}�O��#Jx�p��j0���f����H����6�g~v�ۏ����:�pӫ`���*���U�l�D1�b�x��E�E_�&��<]�=�f�&=1�0���L��Q�d׎�B�&����(�E����H�#�; �<׼�7DZ=zF^�%ѭ��(ps�Cw�gƤ�2����P@�0'�N�Z,x���ٱ�#�_I�Z9)���]�q� �*�OV��ҧl�ԘlFrSvN�(fǴ4E	�+��%��<��� ��b����_�È�]U8� \�^O�V��E����/�3�*h�M��5,#�\��AR1����-���R��T�V��7��fM��V� ����k��r�
Z���򓵅�fq��F��XFt+���w��;�ǎ�N�|%�耱$&�~��RJ�:��&}]������t[�p�(��nks8��D��9�n	�A1���4"�(P:Y)�T�R�Ÿ�����t�	!+E�@��� K0=뾌��#��
Jn�t�����`(�b�MF�R����<!~��%��P���D}�Ңy6�,�o��I��4o�S$45�hN����7�V�H�-1p!�iT0����;ż�w�ϓ�Sd+�3xSl�g�����q��Dfud�NoN�@ď��*��X$�5"a�����$���+Dı+���]����(0ȨiKS^~%�h����#P�_��et�^�2��ޙ�o��_O�EO��#��y��!s�6j�|�9m����-d�uǈJ���GZl����H6�(�;��S�gb$���~�EAV*D� �iC�ݙ�������Q���pK��a;��E�a�ke��o29c�r3z��PP����v�
TЄ��B��V~��}����-(��_iB���0X��j�h��� p�Uj�������EU����tKp��V}T�q�xZ撊���2����T$8Q&(���12���Z�b(�p�~�h��~�~ �lN�h��Xk\�d�#� ��u_�χ���?K&:�d*clZF�=��b&���Jbu��<�񑂥K��J�oa�ʛ�tr�]�g��)W����_��H�%u��{P⼝��������{	"I0K�̠�Tr��>_�t�f���c�����뛵a���{X��a�dga"��&�֔�L�n��0$�ʄC�ӊ�"eW���޴_�]� ��H �g��G��
�Dx����%��C��;�p`2���>�1��lʞQ�)�Gڴe5�2�&�a�
x�n��z>�Uk�(�9�������vMBx�V�i�>K�+tn県EF�טsJĳ����	p[n�/E-��/*Ǜ��������6����H࿂�Hr����B��������(��]���4��`蔍�}���������W�6��5�#z��I��4��g��2����VQݐ���s	�����x��ȧu�W$��g�rx�-@��&E��Wl�g̎��+�I��F�{�Ez5֬���t��7�$�ra��Ƀ�~&��;f��"���/�W��m<DƨR��?+�8�3���}�6=��.��`0J) b� VR�ͳY�K:��x�*�Ŕ�2
���S��H�,*/�}t�(�_ɴVlm=�U�f$�M�'#7�AR�>��N��źq$l�J|���ߌ��x�{�B�cc|d4��ֳJ1W���JE���1!��ά��&��l�E��^
�BD1g�\��{
��Q�Le"�(=���N����g�өJXW��K��s=����TB���qvnOC%��g!��Tk�&qvpL�V�����P����D�;3�	edAc@F۸ ���%�(�������w�
 � �p�&~U΅��Nw)<��d�a(7���\���V�����oR�ҝv�F�b'��ی��.G(ph����y��"�h�;��fY�H5�dU0�R��1W��C�8=wA<G�_�<��r+ӫ�\����6�m�[Ti;K��V/2ƀ���yOv�P72��~�G���^�H�*B>�(;g=B=���T�����[2{;�Rf2P�,w�9�`��I�P%�s����.�l�ǹ#����:cu�i��8ߜN�6/*�K�]��DI'�꠲n����~)w}9� �#��Yx��?�jl�~��;�L󠜷q��p:u�2X��H�*��1��ƪ"̑I�4ѩ�f�q���ݢm�2X�:t"/<rU��b���U�SZ�3�#��`?�5nʈ87�r`���Q�_���?{��HS�(�mp� ��u��#�̏�&���7��3E�0). �����K�_W�&��NO���w/��a��i?P�/���<��9���	��ǭs��_ɕ�	Q��5Y��?��B�,���\?��8g��q�^�sr��������4�S�:E�2N�T��KJE����k9��+MUw:!>X�+;��&���;�˶�(O�
�'��I׮?d�P�^)��N��1�wpf�r�����9ꉅb^ߪ���#r���|
��6qܸ�γ,�_�;��x3�P)�8>_�1���Vjq��Y��<�)%�ojG�6�]7�w�޻s���P�^g
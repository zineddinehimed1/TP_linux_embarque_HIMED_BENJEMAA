��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�/�9�X$+�T�l��h���ɂ����H@� d�}~�A�O����i��q+uC�?���g�-��`��L������xs�>o�}(�Ʈ�l���ٯK�vd�X:6����|<��C��oa�:�P�ؙeV�fp�j�߅�fW�=�M��	:�m����,�t�QE�hY~3�u�ɷ��u�eXJ(�"z3�aG�e��
E�X�X\�M��������j�1���qB'C|�@�$����ϙ��by����S~��>�
�
�Y�
/.��.���k;�6w�{�1RS�P�ϵ�7rʂK�^'K6���[	<'�/��1��ׁ�F[�1p���x�R�.��y�,��u��]�n�KM}��О�&�z�%�4 �,
CEI�=��Jn_h�����*9��&V|��w�7�s�{R2�=�!W#�,�us�<`�Hu.��Q�ɇ��-�Ρ�l抰��N��C� c�K����q�f����Uj�M)�`���;U�i_�B��1~9��y�K�u��i�d�06��\%�� ��=-�dv)'_S=P;�g����y�o��g핉�et��¾�':qWx��W�_LsaJ]��
�=���/��ML��k����}�� �b
��T�UKt;/oY5�?ME��$d6���Z�y(L��&0,UѠ�(�&U\0@���E�`��7ɫ��F~
KP2dd�5'ou�jX,�z{I��q���=�V���Mq�d}���4Tں�KÃpQ��׊����Q|vMnTU�Q�� u|r��8]������* ��Lٺk�ʅ+,��5a�r7p���p�&�6��<���LqF��X���+�Tr���+FMY�{�Z�����9X�S툱�@
�����
��2��D��A����M�Ǳ���`�!�?���1�u�a;��lt���A�<I�?�$I�_ԟ�X�l�����ڵ��@��zX1\AA��=z��C��+\i�����M�q��ݚ��Ӯ��K�������M/o���J< 뒵,xO��������������m�s�/�\�Ҧ�����lPO?�bZ=���J2)� ��F��E�9��%]�к(zn�XF]b��Iy2z{�S��D:�@k!��̷�c�1M�1.2X���|X�4S��~�m�w���r�ߪ�����V_ֶ�����0��7J7�ޫ|�%Q>O�	H���B��&$ۿ�[!�@�����w���l��2`�`l����6��Z=�& -!d'�#!�0������ǠXϷN}/���ǤYqC��_�8�*�Q ���n��g���&��}/���R�,��i^B
v�Xx���=�.�y� ;��W�3�X{\6��1s5�,��D8x�$ ��:E"O����ߗ��	�nI�v:!d�JD
8�c1��e�-n���c_��]��